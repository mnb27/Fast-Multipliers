`timescale 1ns / 1ps

module GenPPRow0(x,y,a0b0,a1b0,a2b0,a3b0,a4b0,a5b0,a6b0,a7b0,a8b0,a9b0,a10b0,a11b0,a12b0,a13b0,a14b0,a15b0,a16b0,a17b0,a18b0,a19b0,a20b0,a21b0,a22b0,a23b0,a24b0,a25b0,a26b0,a27b0,a28b0,a29b0,a30b0,a31b0);
input [31:0] x;
input y;
output reg a0b0,a1b0,a2b0,a3b0,a4b0,a5b0,a6b0,a7b0,a8b0,a9b0,a10b0,a11b0,a12b0,a13b0,a14b0,a15b0,a16b0,a17b0,a18b0,a19b0,a20b0,a21b0,a22b0,a23b0,a24b0,a25b0,a26b0,a27b0,a28b0,a29b0,a30b0,a31b0;

always@(x,y)begin
	a0b0 <= x[0] & y;
	a1b0 <= x[1] & y;
	a2b0 <= x[2] & y;
	a3b0 <= x[3] & y;
	a4b0 <= x[4] & y;
	a5b0 <= x[5] & y;
	a6b0 <= x[6] & y;
	a7b0 <= x[7] & y;
	a8b0 <= x[8] & y;
	a9b0 <= x[9] & y;
	a10b0 <= x[10] & y;
	a11b0 <= x[11] & y;
	a12b0 <= x[12] & y;
	a13b0 <= x[13] & y;
	a14b0 <= x[14] & y;
	a15b0 <= x[15] & y;
	a16b0 <= x[16] & y;
	a17b0 <= x[17] & y;
	a18b0 <= x[18] & y;
	a19b0 <= x[19] & y;
	a20b0 <= x[20] & y;
	a21b0 <= x[21] & y;
	a22b0 <= x[22] & y;
	a23b0 <= x[23] & y;
	a24b0 <= x[24] & y;
	a25b0 <= x[25] & y;
	a26b0 <= x[26] & y;
	a27b0 <= x[27] & y;
	a28b0 <= x[28] & y;
	a29b0 <= x[29] & y;
	a30b0 <= x[30] & y;
	a31b0 <= x[31] & y;
end

endmodule

module GenPPRow1(x,y,a0b1,a1b1,a2b1,a3b1,a4b1,a5b1,a6b1,a7b1,a8b1,a9b1,a10b1,a11b1,a12b1,a13b1,a14b1,a15b1,a16b1,a17b1,a18b1,a19b1,a20b1,a21b1,a22b1,a23b1,a24b1,a25b1,a26b1,a27b1,a28b1,a29b1,a30b1,a31b1);
input [31:0] x;
input y;
output reg a0b1,a1b1,a2b1,a3b1,a4b1,a5b1,a6b1,a7b1,a8b1,a9b1,a10b1,a11b1,a12b1,a13b1,a14b1,a15b1,a16b1,a17b1,a18b1,a19b1,a20b1,a21b1,a22b1,a23b1,a24b1,a25b1,a26b1,a27b1,a28b1,a29b1,a30b1,a31b1;

always@(x,y)begin
	a0b1 <= x[0] & y;
	a1b1 <= x[1] & y;
	a2b1 <= x[2] & y;
	a3b1 <= x[3] & y;
	a4b1 <= x[4] & y;
	a5b1 <= x[5] & y;
	a6b1 <= x[6] & y;
	a7b1 <= x[7] & y;
	a8b1 <= x[8] & y;
	a9b1 <= x[9] & y;
	a10b1 <= x[10] & y;
	a11b1 <= x[11] & y;
	a12b1 <= x[12] & y;
	a13b1 <= x[13] & y;
	a14b1 <= x[14] & y;
	a15b1 <= x[15] & y;
	a16b1 <= x[16] & y;
	a17b1 <= x[17] & y;
	a18b1 <= x[18] & y;
	a19b1 <= x[19] & y;
	a20b1 <= x[20] & y;
	a21b1 <= x[21] & y;
	a22b1 <= x[22] & y;
	a23b1 <= x[23] & y;
	a24b1 <= x[24] & y;
	a25b1 <= x[25] & y;
	a26b1 <= x[26] & y;
	a27b1 <= x[27] & y;
	a28b1 <= x[28] & y;
	a29b1 <= x[29] & y;
	a30b1 <= x[30] & y;
	a31b1 <= x[31] & y;
end

endmodule

module GenPPRow2(x,y,a0b2,a1b2,a2b2,a3b2,a4b2,a5b2,a6b2,a7b2,a8b2,a9b2,a10b2,a11b2,a12b2,a13b2,a14b2,a15b2,a16b2,a17b2,a18b2,a19b2,a20b2,a21b2,a22b2,a23b2,a24b2,a25b2,a26b2,a27b2,a28b2,a29b2,a30b2,a31b2);
input [31:0] x;
input y;
output reg a0b2,a1b2,a2b2,a3b2,a4b2,a5b2,a6b2,a7b2,a8b2,a9b2,a10b2,a11b2,a12b2,a13b2,a14b2,a15b2,a16b2,a17b2,a18b2,a19b2,a20b2,a21b2,a22b2,a23b2,a24b2,a25b2,a26b2,a27b2,a28b2,a29b2,a30b2,a31b2;

always@(x,y)begin
	a0b2 <= x[0] & y;
	a1b2 <= x[1] & y;
	a2b2 <= x[2] & y;
	a3b2 <= x[3] & y;
	a4b2 <= x[4] & y;
	a5b2 <= x[5] & y;
	a6b2 <= x[6] & y;
	a7b2 <= x[7] & y;
	a8b2 <= x[8] & y;
	a9b2 <= x[9] & y;
	a10b2 <= x[10] & y;
	a11b2 <= x[11] & y;
	a12b2 <= x[12] & y;
	a13b2 <= x[13] & y;
	a14b2 <= x[14] & y;
	a15b2 <= x[15] & y;
	a16b2 <= x[16] & y;
	a17b2 <= x[17] & y;
	a18b2 <= x[18] & y;
	a19b2 <= x[19] & y;
	a20b2 <= x[20] & y;
	a21b2 <= x[21] & y;
	a22b2 <= x[22] & y;
	a23b2 <= x[23] & y;
	a24b2 <= x[24] & y;
	a25b2 <= x[25] & y;
	a26b2 <= x[26] & y;
	a27b2 <= x[27] & y;
	a28b2 <= x[28] & y;
	a29b2 <= x[29] & y;
	a30b2 <= x[30] & y;
	a31b2 <= x[31] & y;
end

endmodule

module GenPPRow3(x,y,a0b3,a1b3,a2b3,a3b3,a4b3,a5b3,a6b3,a7b3,a8b3,a9b3,a10b3,a11b3,a12b3,a13b3,a14b3,a15b3,a16b3,a17b3,a18b3,a19b3,a20b3,a21b3,a22b3,a23b3,a24b3,a25b3,a26b3,a27b3,a28b3,a29b3,a30b3,a31b3);
input [31:0] x;
input y;
output reg a0b3,a1b3,a2b3,a3b3,a4b3,a5b3,a6b3,a7b3,a8b3,a9b3,a10b3,a11b3,a12b3,a13b3,a14b3,a15b3,a16b3,a17b3,a18b3,a19b3,a20b3,a21b3,a22b3,a23b3,a24b3,a25b3,a26b3,a27b3,a28b3,a29b3,a30b3,a31b3;

always@(x,y)begin
	a0b3 <= x[0] & y;
	a1b3 <= x[1] & y;
	a2b3 <= x[2] & y;
	a3b3 <= x[3] & y;
	a4b3 <= x[4] & y;
	a5b3 <= x[5] & y;
	a6b3 <= x[6] & y;
	a7b3 <= x[7] & y;
	a8b3 <= x[8] & y;
	a9b3 <= x[9] & y;
	a10b3 <= x[10] & y;
	a11b3 <= x[11] & y;
	a12b3 <= x[12] & y;
	a13b3 <= x[13] & y;
	a14b3 <= x[14] & y;
	a15b3 <= x[15] & y;
	a16b3 <= x[16] & y;
	a17b3 <= x[17] & y;
	a18b3 <= x[18] & y;
	a19b3 <= x[19] & y;
	a20b3 <= x[20] & y;
	a21b3 <= x[21] & y;
	a22b3 <= x[22] & y;
	a23b3 <= x[23] & y;
	a24b3 <= x[24] & y;
	a25b3 <= x[25] & y;
	a26b3 <= x[26] & y;
	a27b3 <= x[27] & y;
	a28b3 <= x[28] & y;
	a29b3 <= x[29] & y;
	a30b3 <= x[30] & y;
	a31b3 <= x[31] & y;
end

endmodule

module GenPPRow4(x,y,a0b4,a1b4,a2b4,a3b4,a4b4,a5b4,a6b4,a7b4,a8b4,a9b4,a10b4,a11b4,a12b4,a13b4,a14b4,a15b4,a16b4,a17b4,a18b4,a19b4,a20b4,a21b4,a22b4,a23b4,a24b4,a25b4,a26b4,a27b4,a28b4,a29b4,a30b4,a31b4);
input [31:0] x;
input y;
output reg a0b4,a1b4,a2b4,a3b4,a4b4,a5b4,a6b4,a7b4,a8b4,a9b4,a10b4,a11b4,a12b4,a13b4,a14b4,a15b4,a16b4,a17b4,a18b4,a19b4,a20b4,a21b4,a22b4,a23b4,a24b4,a25b4,a26b4,a27b4,a28b4,a29b4,a30b4,a31b4;

always@(x,y)begin
	a0b4 <= x[0] & y;
	a1b4 <= x[1] & y;
	a2b4 <= x[2] & y;
	a3b4 <= x[3] & y;
	a4b4 <= x[4] & y;
	a5b4 <= x[5] & y;
	a6b4 <= x[6] & y;
	a7b4 <= x[7] & y;
	a8b4 <= x[8] & y;
	a9b4 <= x[9] & y;
	a10b4 <= x[10] & y;
	a11b4 <= x[11] & y;
	a12b4 <= x[12] & y;
	a13b4 <= x[13] & y;
	a14b4 <= x[14] & y;
	a15b4 <= x[15] & y;
	a16b4 <= x[16] & y;
	a17b4 <= x[17] & y;
	a18b4 <= x[18] & y;
	a19b4 <= x[19] & y;
	a20b4 <= x[20] & y;
	a21b4 <= x[21] & y;
	a22b4 <= x[22] & y;
	a23b4 <= x[23] & y;
	a24b4 <= x[24] & y;
	a25b4 <= x[25] & y;
	a26b4 <= x[26] & y;
	a27b4 <= x[27] & y;
	a28b4 <= x[28] & y;
	a29b4 <= x[29] & y;
	a30b4 <= x[30] & y;
	a31b4 <= x[31] & y;
end

endmodule

module GenPPRow5(x,y,a0b5,a1b5,a2b5,a3b5,a4b5,a5b5,a6b5,a7b5,a8b5,a9b5,a10b5,a11b5,a12b5,a13b5,a14b5,a15b5,a16b5,a17b5,a18b5,a19b5,a20b5,a21b5,a22b5,a23b5,a24b5,a25b5,a26b5,a27b5,a28b5,a29b5,a30b5,a31b5);
input [31:0] x;
input y;
output reg a0b5,a1b5,a2b5,a3b5,a4b5,a5b5,a6b5,a7b5,a8b5,a9b5,a10b5,a11b5,a12b5,a13b5,a14b5,a15b5,a16b5,a17b5,a18b5,a19b5,a20b5,a21b5,a22b5,a23b5,a24b5,a25b5,a26b5,a27b5,a28b5,a29b5,a30b5,a31b5;

always@(x,y)begin
	a0b5 <= x[0] & y;
	a1b5 <= x[1] & y;
	a2b5 <= x[2] & y;
	a3b5 <= x[3] & y;
	a4b5 <= x[4] & y;
	a5b5 <= x[5] & y;
	a6b5 <= x[6] & y;
	a7b5 <= x[7] & y;
	a8b5 <= x[8] & y;
	a9b5 <= x[9] & y;
	a10b5 <= x[10] & y;
	a11b5 <= x[11] & y;
	a12b5 <= x[12] & y;
	a13b5 <= x[13] & y;
	a14b5 <= x[14] & y;
	a15b5 <= x[15] & y;
	a16b5 <= x[16] & y;
	a17b5 <= x[17] & y;
	a18b5 <= x[18] & y;
	a19b5 <= x[19] & y;
	a20b5 <= x[20] & y;
	a21b5 <= x[21] & y;
	a22b5 <= x[22] & y;
	a23b5 <= x[23] & y;
	a24b5 <= x[24] & y;
	a25b5 <= x[25] & y;
	a26b5 <= x[26] & y;
	a27b5 <= x[27] & y;
	a28b5 <= x[28] & y;
	a29b5 <= x[29] & y;
	a30b5 <= x[30] & y;
	a31b5 <= x[31] & y;
end

endmodule

module GenPPRow6(x,y,a0b6,a1b6,a2b6,a3b6,a4b6,a5b6,a6b6,a7b6,a8b6,a9b6,a10b6,a11b6,a12b6,a13b6,a14b6,a15b6,a16b6,a17b6,a18b6,a19b6,a20b6,a21b6,a22b6,a23b6,a24b6,a25b6,a26b6,a27b6,a28b6,a29b6,a30b6,a31b6);
input [31:0] x;
input y;
output reg a0b6,a1b6,a2b6,a3b6,a4b6,a5b6,a6b6,a7b6,a8b6,a9b6,a10b6,a11b6,a12b6,a13b6,a14b6,a15b6,a16b6,a17b6,a18b6,a19b6,a20b6,a21b6,a22b6,a23b6,a24b6,a25b6,a26b6,a27b6,a28b6,a29b6,a30b6,a31b6;

always@(x,y)begin
	a0b6 <= x[0] & y;
	a1b6 <= x[1] & y;
	a2b6 <= x[2] & y;
	a3b6 <= x[3] & y;
	a4b6 <= x[4] & y;
	a5b6 <= x[5] & y;
	a6b6 <= x[6] & y;
	a7b6 <= x[7] & y;
	a8b6 <= x[8] & y;
	a9b6 <= x[9] & y;
	a10b6 <= x[10] & y;
	a11b6 <= x[11] & y;
	a12b6 <= x[12] & y;
	a13b6 <= x[13] & y;
	a14b6 <= x[14] & y;
	a15b6 <= x[15] & y;
	a16b6 <= x[16] & y;
	a17b6 <= x[17] & y;
	a18b6 <= x[18] & y;
	a19b6 <= x[19] & y;
	a20b6 <= x[20] & y;
	a21b6 <= x[21] & y;
	a22b6 <= x[22] & y;
	a23b6 <= x[23] & y;
	a24b6 <= x[24] & y;
	a25b6 <= x[25] & y;
	a26b6 <= x[26] & y;
	a27b6 <= x[27] & y;
	a28b6 <= x[28] & y;
	a29b6 <= x[29] & y;
	a30b6 <= x[30] & y;
	a31b6 <= x[31] & y;
end

endmodule

module GenPPRow7(x,y,a0b7,a1b7,a2b7,a3b7,a4b7,a5b7,a6b7,a7b7,a8b7,a9b7,a10b7,a11b7,a12b7,a13b7,a14b7,a15b7,a16b7,a17b7,a18b7,a19b7,a20b7,a21b7,a22b7,a23b7,a24b7,a25b7,a26b7,a27b7,a28b7,a29b7,a30b7,a31b7);
input [31:0] x;
input y;
output reg a0b7,a1b7,a2b7,a3b7,a4b7,a5b7,a6b7,a7b7,a8b7,a9b7,a10b7,a11b7,a12b7,a13b7,a14b7,a15b7,a16b7,a17b7,a18b7,a19b7,a20b7,a21b7,a22b7,a23b7,a24b7,a25b7,a26b7,a27b7,a28b7,a29b7,a30b7,a31b7;

always@(x,y)begin
	a0b7 <= x[0] & y;
	a1b7 <= x[1] & y;
	a2b7 <= x[2] & y;
	a3b7 <= x[3] & y;
	a4b7 <= x[4] & y;
	a5b7 <= x[5] & y;
	a6b7 <= x[6] & y;
	a7b7 <= x[7] & y;
	a8b7 <= x[8] & y;
	a9b7 <= x[9] & y;
	a10b7 <= x[10] & y;
	a11b7 <= x[11] & y;
	a12b7 <= x[12] & y;
	a13b7 <= x[13] & y;
	a14b7 <= x[14] & y;
	a15b7 <= x[15] & y;
	a16b7 <= x[16] & y;
	a17b7 <= x[17] & y;
	a18b7 <= x[18] & y;
	a19b7 <= x[19] & y;
	a20b7 <= x[20] & y;
	a21b7 <= x[21] & y;
	a22b7 <= x[22] & y;
	a23b7 <= x[23] & y;
	a24b7 <= x[24] & y;
	a25b7 <= x[25] & y;
	a26b7 <= x[26] & y;
	a27b7 <= x[27] & y;
	a28b7 <= x[28] & y;
	a29b7 <= x[29] & y;
	a30b7 <= x[30] & y;
	a31b7 <= x[31] & y;
end

endmodule

module GenPPRow8(x,y,a0b8,a1b8,a2b8,a3b8,a4b8,a5b8,a6b8,a7b8,a8b8,a9b8,a10b8,a11b8,a12b8,a13b8,a14b8,a15b8,a16b8,a17b8,a18b8,a19b8,a20b8,a21b8,a22b8,a23b8,a24b8,a25b8,a26b8,a27b8,a28b8,a29b8,a30b8,a31b8);
input [31:0] x;
input y;
output reg a0b8,a1b8,a2b8,a3b8,a4b8,a5b8,a6b8,a7b8,a8b8,a9b8,a10b8,a11b8,a12b8,a13b8,a14b8,a15b8,a16b8,a17b8,a18b8,a19b8,a20b8,a21b8,a22b8,a23b8,a24b8,a25b8,a26b8,a27b8,a28b8,a29b8,a30b8,a31b8;

always@(x,y)begin
	a0b8 <= x[0] & y;
	a1b8 <= x[1] & y;
	a2b8 <= x[2] & y;
	a3b8 <= x[3] & y;
	a4b8 <= x[4] & y;
	a5b8 <= x[5] & y;
	a6b8 <= x[6] & y;
	a7b8 <= x[7] & y;
	a8b8 <= x[8] & y;
	a9b8 <= x[9] & y;
	a10b8 <= x[10] & y;
	a11b8 <= x[11] & y;
	a12b8 <= x[12] & y;
	a13b8 <= x[13] & y;
	a14b8 <= x[14] & y;
	a15b8 <= x[15] & y;
	a16b8 <= x[16] & y;
	a17b8 <= x[17] & y;
	a18b8 <= x[18] & y;
	a19b8 <= x[19] & y;
	a20b8 <= x[20] & y;
	a21b8 <= x[21] & y;
	a22b8 <= x[22] & y;
	a23b8 <= x[23] & y;
	a24b8 <= x[24] & y;
	a25b8 <= x[25] & y;
	a26b8 <= x[26] & y;
	a27b8 <= x[27] & y;
	a28b8 <= x[28] & y;
	a29b8 <= x[29] & y;
	a30b8 <= x[30] & y;
	a31b8 <= x[31] & y;
end

endmodule

module GenPPRow9(x,y,a0b9,a1b9,a2b9,a3b9,a4b9,a5b9,a6b9,a7b9,a8b9,a9b9,a10b9,a11b9,a12b9,a13b9,a14b9,a15b9,a16b9,a17b9,a18b9,a19b9,a20b9,a21b9,a22b9,a23b9,a24b9,a25b9,a26b9,a27b9,a28b9,a29b9,a30b9,a31b9);
input [31:0] x;
input y;
output reg a0b9,a1b9,a2b9,a3b9,a4b9,a5b9,a6b9,a7b9,a8b9,a9b9,a10b9,a11b9,a12b9,a13b9,a14b9,a15b9,a16b9,a17b9,a18b9,a19b9,a20b9,a21b9,a22b9,a23b9,a24b9,a25b9,a26b9,a27b9,a28b9,a29b9,a30b9,a31b9;

always@(x,y)begin
	a0b9 <= x[0] & y;
	a1b9 <= x[1] & y;
	a2b9 <= x[2] & y;
	a3b9 <= x[3] & y;
	a4b9 <= x[4] & y;
	a5b9 <= x[5] & y;
	a6b9 <= x[6] & y;
	a7b9 <= x[7] & y;
	a8b9 <= x[8] & y;
	a9b9 <= x[9] & y;
	a10b9 <= x[10] & y;
	a11b9 <= x[11] & y;
	a12b9 <= x[12] & y;
	a13b9 <= x[13] & y;
	a14b9 <= x[14] & y;
	a15b9 <= x[15] & y;
	a16b9 <= x[16] & y;
	a17b9 <= x[17] & y;
	a18b9 <= x[18] & y;
	a19b9 <= x[19] & y;
	a20b9 <= x[20] & y;
	a21b9 <= x[21] & y;
	a22b9 <= x[22] & y;
	a23b9 <= x[23] & y;
	a24b9 <= x[24] & y;
	a25b9 <= x[25] & y;
	a26b9 <= x[26] & y;
	a27b9 <= x[27] & y;
	a28b9 <= x[28] & y;
	a29b9 <= x[29] & y;
	a30b9 <= x[30] & y;
	a31b9 <= x[31] & y;
end

endmodule

module GenPPRow10(x,y,a0b10,a1b10,a2b10,a3b10,a4b10,a5b10,a6b10,a7b10,a8b10,a9b10,a10b10,a11b10,a12b10,a13b10,a14b10,a15b10,a16b10,a17b10,a18b10,a19b10,a20b10,a21b10,a22b10,a23b10,a24b10,a25b10,a26b10,a27b10,a28b10,a29b10,a30b10,a31b10);
input [31:0] x;
input y;
output reg a0b10,a1b10,a2b10,a3b10,a4b10,a5b10,a6b10,a7b10,a8b10,a9b10,a10b10,a11b10,a12b10,a13b10,a14b10,a15b10,a16b10,a17b10,a18b10,a19b10,a20b10,a21b10,a22b10,a23b10,a24b10,a25b10,a26b10,a27b10,a28b10,a29b10,a30b10,a31b10;

always@(x,y)begin
	a0b10 <= x[0] & y;
	a1b10 <= x[1] & y;
	a2b10 <= x[2] & y;
	a3b10 <= x[3] & y;
	a4b10 <= x[4] & y;
	a5b10 <= x[5] & y;
	a6b10 <= x[6] & y;
	a7b10 <= x[7] & y;
	a8b10 <= x[8] & y;
	a9b10 <= x[9] & y;
	a10b10 <= x[10] & y;
	a11b10 <= x[11] & y;
	a12b10 <= x[12] & y;
	a13b10 <= x[13] & y;
	a14b10 <= x[14] & y;
	a15b10 <= x[15] & y;
	a16b10 <= x[16] & y;
	a17b10 <= x[17] & y;
	a18b10 <= x[18] & y;
	a19b10 <= x[19] & y;
	a20b10 <= x[20] & y;
	a21b10 <= x[21] & y;
	a22b10 <= x[22] & y;
	a23b10 <= x[23] & y;
	a24b10 <= x[24] & y;
	a25b10 <= x[25] & y;
	a26b10 <= x[26] & y;
	a27b10 <= x[27] & y;
	a28b10 <= x[28] & y;
	a29b10 <= x[29] & y;
	a30b10 <= x[30] & y;
	a31b10 <= x[31] & y;
end

endmodule

module GenPPRow11(x,y,a0b11,a1b11,a2b11,a3b11,a4b11,a5b11,a6b11,a7b11,a8b11,a9b11,a10b11,a11b11,a12b11,a13b11,a14b11,a15b11,a16b11,a17b11,a18b11,a19b11,a20b11,a21b11,a22b11,a23b11,a24b11,a25b11,a26b11,a27b11,a28b11,a29b11,a30b11,a31b11);
input [31:0] x;
input y;
output reg a0b11,a1b11,a2b11,a3b11,a4b11,a5b11,a6b11,a7b11,a8b11,a9b11,a10b11,a11b11,a12b11,a13b11,a14b11,a15b11,a16b11,a17b11,a18b11,a19b11,a20b11,a21b11,a22b11,a23b11,a24b11,a25b11,a26b11,a27b11,a28b11,a29b11,a30b11,a31b11;

always@(x,y)begin
	a0b11 <= x[0] & y;
	a1b11 <= x[1] & y;
	a2b11 <= x[2] & y;
	a3b11 <= x[3] & y;
	a4b11 <= x[4] & y;
	a5b11 <= x[5] & y;
	a6b11 <= x[6] & y;
	a7b11 <= x[7] & y;
	a8b11 <= x[8] & y;
	a9b11 <= x[9] & y;
	a10b11 <= x[10] & y;
	a11b11 <= x[11] & y;
	a12b11 <= x[12] & y;
	a13b11 <= x[13] & y;
	a14b11 <= x[14] & y;
	a15b11 <= x[15] & y;
	a16b11 <= x[16] & y;
	a17b11 <= x[17] & y;
	a18b11 <= x[18] & y;
	a19b11 <= x[19] & y;
	a20b11 <= x[20] & y;
	a21b11 <= x[21] & y;
	a22b11 <= x[22] & y;
	a23b11 <= x[23] & y;
	a24b11 <= x[24] & y;
	a25b11 <= x[25] & y;
	a26b11 <= x[26] & y;
	a27b11 <= x[27] & y;
	a28b11 <= x[28] & y;
	a29b11 <= x[29] & y;
	a30b11 <= x[30] & y;
	a31b11 <= x[31] & y;
end

endmodule

module GenPPRow12(x,y,a0b12,a1b12,a2b12,a3b12,a4b12,a5b12,a6b12,a7b12,a8b12,a9b12,a10b12,a11b12,a12b12,a13b12,a14b12,a15b12,a16b12,a17b12,a18b12,a19b12,a20b12,a21b12,a22b12,a23b12,a24b12,a25b12,a26b12,a27b12,a28b12,a29b12,a30b12,a31b12);
input [31:0] x;
input y;
output reg a0b12,a1b12,a2b12,a3b12,a4b12,a5b12,a6b12,a7b12,a8b12,a9b12,a10b12,a11b12,a12b12,a13b12,a14b12,a15b12,a16b12,a17b12,a18b12,a19b12,a20b12,a21b12,a22b12,a23b12,a24b12,a25b12,a26b12,a27b12,a28b12,a29b12,a30b12,a31b12;

always@(x,y)begin
	a0b12 <= x[0] & y;
	a1b12 <= x[1] & y;
	a2b12 <= x[2] & y;
	a3b12 <= x[3] & y;
	a4b12 <= x[4] & y;
	a5b12 <= x[5] & y;
	a6b12 <= x[6] & y;
	a7b12 <= x[7] & y;
	a8b12 <= x[8] & y;
	a9b12 <= x[9] & y;
	a10b12 <= x[10] & y;
	a11b12 <= x[11] & y;
	a12b12 <= x[12] & y;
	a13b12 <= x[13] & y;
	a14b12 <= x[14] & y;
	a15b12 <= x[15] & y;
	a16b12 <= x[16] & y;
	a17b12 <= x[17] & y;
	a18b12 <= x[18] & y;
	a19b12 <= x[19] & y;
	a20b12 <= x[20] & y;
	a21b12 <= x[21] & y;
	a22b12 <= x[22] & y;
	a23b12 <= x[23] & y;
	a24b12 <= x[24] & y;
	a25b12 <= x[25] & y;
	a26b12 <= x[26] & y;
	a27b12 <= x[27] & y;
	a28b12 <= x[28] & y;
	a29b12 <= x[29] & y;
	a30b12 <= x[30] & y;
	a31b12 <= x[31] & y;
end

endmodule

module GenPPRow13(x,y,a0b13,a1b13,a2b13,a3b13,a4b13,a5b13,a6b13,a7b13,a8b13,a9b13,a10b13,a11b13,a12b13,a13b13,a14b13,a15b13,a16b13,a17b13,a18b13,a19b13,a20b13,a21b13,a22b13,a23b13,a24b13,a25b13,a26b13,a27b13,a28b13,a29b13,a30b13,a31b13);
input [31:0] x;
input y;
output reg a0b13,a1b13,a2b13,a3b13,a4b13,a5b13,a6b13,a7b13,a8b13,a9b13,a10b13,a11b13,a12b13,a13b13,a14b13,a15b13,a16b13,a17b13,a18b13,a19b13,a20b13,a21b13,a22b13,a23b13,a24b13,a25b13,a26b13,a27b13,a28b13,a29b13,a30b13,a31b13;

always@(x,y)begin
	a0b13 <= x[0] & y;
	a1b13 <= x[1] & y;
	a2b13 <= x[2] & y;
	a3b13 <= x[3] & y;
	a4b13 <= x[4] & y;
	a5b13 <= x[5] & y;
	a6b13 <= x[6] & y;
	a7b13 <= x[7] & y;
	a8b13 <= x[8] & y;
	a9b13 <= x[9] & y;
	a10b13 <= x[10] & y;
	a11b13 <= x[11] & y;
	a12b13 <= x[12] & y;
	a13b13 <= x[13] & y;
	a14b13 <= x[14] & y;
	a15b13 <= x[15] & y;
	a16b13 <= x[16] & y;
	a17b13 <= x[17] & y;
	a18b13 <= x[18] & y;
	a19b13 <= x[19] & y;
	a20b13 <= x[20] & y;
	a21b13 <= x[21] & y;
	a22b13 <= x[22] & y;
	a23b13 <= x[23] & y;
	a24b13 <= x[24] & y;
	a25b13 <= x[25] & y;
	a26b13 <= x[26] & y;
	a27b13 <= x[27] & y;
	a28b13 <= x[28] & y;
	a29b13 <= x[29] & y;
	a30b13 <= x[30] & y;
	a31b13 <= x[31] & y;
end

endmodule

module GenPPRow14(x,y,a0b14,a1b14,a2b14,a3b14,a4b14,a5b14,a6b14,a7b14,a8b14,a9b14,a10b14,a11b14,a12b14,a13b14,a14b14,a15b14,a16b14,a17b14,a18b14,a19b14,a20b14,a21b14,a22b14,a23b14,a24b14,a25b14,a26b14,a27b14,a28b14,a29b14,a30b14,a31b14);
input [31:0] x;
input y;
output reg a0b14,a1b14,a2b14,a3b14,a4b14,a5b14,a6b14,a7b14,a8b14,a9b14,a10b14,a11b14,a12b14,a13b14,a14b14,a15b14,a16b14,a17b14,a18b14,a19b14,a20b14,a21b14,a22b14,a23b14,a24b14,a25b14,a26b14,a27b14,a28b14,a29b14,a30b14,a31b14;

always@(x,y)begin
	a0b14 <= x[0] & y;
	a1b14 <= x[1] & y;
	a2b14 <= x[2] & y;
	a3b14 <= x[3] & y;
	a4b14 <= x[4] & y;
	a5b14 <= x[5] & y;
	a6b14 <= x[6] & y;
	a7b14 <= x[7] & y;
	a8b14 <= x[8] & y;
	a9b14 <= x[9] & y;
	a10b14 <= x[10] & y;
	a11b14 <= x[11] & y;
	a12b14 <= x[12] & y;
	a13b14 <= x[13] & y;
	a14b14 <= x[14] & y;
	a15b14 <= x[15] & y;
	a16b14 <= x[16] & y;
	a17b14 <= x[17] & y;
	a18b14 <= x[18] & y;
	a19b14 <= x[19] & y;
	a20b14 <= x[20] & y;
	a21b14 <= x[21] & y;
	a22b14 <= x[22] & y;
	a23b14 <= x[23] & y;
	a24b14 <= x[24] & y;
	a25b14 <= x[25] & y;
	a26b14 <= x[26] & y;
	a27b14 <= x[27] & y;
	a28b14 <= x[28] & y;
	a29b14 <= x[29] & y;
	a30b14 <= x[30] & y;
	a31b14 <= x[31] & y;
end

endmodule

module GenPPRow15(x,y,a0b15,a1b15,a2b15,a3b15,a4b15,a5b15,a6b15,a7b15,a8b15,a9b15,a10b15,a11b15,a12b15,a13b15,a14b15,a15b15,a16b15,a17b15,a18b15,a19b15,a20b15,a21b15,a22b15,a23b15,a24b15,a25b15,a26b15,a27b15,a28b15,a29b15,a30b15,a31b15);
input [31:0] x;
input y;
output reg a0b15,a1b15,a2b15,a3b15,a4b15,a5b15,a6b15,a7b15,a8b15,a9b15,a10b15,a11b15,a12b15,a13b15,a14b15,a15b15,a16b15,a17b15,a18b15,a19b15,a20b15,a21b15,a22b15,a23b15,a24b15,a25b15,a26b15,a27b15,a28b15,a29b15,a30b15,a31b15;

always@(x,y)begin
	a0b15 <= x[0] & y;
	a1b15 <= x[1] & y;
	a2b15 <= x[2] & y;
	a3b15 <= x[3] & y;
	a4b15 <= x[4] & y;
	a5b15 <= x[5] & y;
	a6b15 <= x[6] & y;
	a7b15 <= x[7] & y;
	a8b15 <= x[8] & y;
	a9b15 <= x[9] & y;
	a10b15 <= x[10] & y;
	a11b15 <= x[11] & y;
	a12b15 <= x[12] & y;
	a13b15 <= x[13] & y;
	a14b15 <= x[14] & y;
	a15b15 <= x[15] & y;
	a16b15 <= x[16] & y;
	a17b15 <= x[17] & y;
	a18b15 <= x[18] & y;
	a19b15 <= x[19] & y;
	a20b15 <= x[20] & y;
	a21b15 <= x[21] & y;
	a22b15 <= x[22] & y;
	a23b15 <= x[23] & y;
	a24b15 <= x[24] & y;
	a25b15 <= x[25] & y;
	a26b15 <= x[26] & y;
	a27b15 <= x[27] & y;
	a28b15 <= x[28] & y;
	a29b15 <= x[29] & y;
	a30b15 <= x[30] & y;
	a31b15 <= x[31] & y;
end

endmodule

module GenPPRow16(x,y,a0b16,a1b16,a2b16,a3b16,a4b16,a5b16,a6b16,a7b16,a8b16,a9b16,a10b16,a11b16,a12b16,a13b16,a14b16,a15b16,a16b16,a17b16,a18b16,a19b16,a20b16,a21b16,a22b16,a23b16,a24b16,a25b16,a26b16,a27b16,a28b16,a29b16,a30b16,a31b16);
input [31:0] x;
input y;
output reg a0b16,a1b16,a2b16,a3b16,a4b16,a5b16,a6b16,a7b16,a8b16,a9b16,a10b16,a11b16,a12b16,a13b16,a14b16,a15b16,a16b16,a17b16,a18b16,a19b16,a20b16,a21b16,a22b16,a23b16,a24b16,a25b16,a26b16,a27b16,a28b16,a29b16,a30b16,a31b16;

always@(x,y)begin
	a0b16 <= x[0] & y;
	a1b16 <= x[1] & y;
	a2b16 <= x[2] & y;
	a3b16 <= x[3] & y;
	a4b16 <= x[4] & y;
	a5b16 <= x[5] & y;
	a6b16 <= x[6] & y;
	a7b16 <= x[7] & y;
	a8b16 <= x[8] & y;
	a9b16 <= x[9] & y;
	a10b16 <= x[10] & y;
	a11b16 <= x[11] & y;
	a12b16 <= x[12] & y;
	a13b16 <= x[13] & y;
	a14b16 <= x[14] & y;
	a15b16 <= x[15] & y;
	a16b16 <= x[16] & y;
	a17b16 <= x[17] & y;
	a18b16 <= x[18] & y;
	a19b16 <= x[19] & y;
	a20b16 <= x[20] & y;
	a21b16 <= x[21] & y;
	a22b16 <= x[22] & y;
	a23b16 <= x[23] & y;
	a24b16 <= x[24] & y;
	a25b16 <= x[25] & y;
	a26b16 <= x[26] & y;
	a27b16 <= x[27] & y;
	a28b16 <= x[28] & y;
	a29b16 <= x[29] & y;
	a30b16 <= x[30] & y;
	a31b16 <= x[31] & y;
end

endmodule

module GenPPRow17(x,y,a0b17,a1b17,a2b17,a3b17,a4b17,a5b17,a6b17,a7b17,a8b17,a9b17,a10b17,a11b17,a12b17,a13b17,a14b17,a15b17,a16b17,a17b17,a18b17,a19b17,a20b17,a21b17,a22b17,a23b17,a24b17,a25b17,a26b17,a27b17,a28b17,a29b17,a30b17,a31b17);
input [31:0] x;
input y;
output reg a0b17,a1b17,a2b17,a3b17,a4b17,a5b17,a6b17,a7b17,a8b17,a9b17,a10b17,a11b17,a12b17,a13b17,a14b17,a15b17,a16b17,a17b17,a18b17,a19b17,a20b17,a21b17,a22b17,a23b17,a24b17,a25b17,a26b17,a27b17,a28b17,a29b17,a30b17,a31b17;

always@(x,y)begin
	a0b17 <= x[0] & y;
	a1b17 <= x[1] & y;
	a2b17 <= x[2] & y;
	a3b17 <= x[3] & y;
	a4b17 <= x[4] & y;
	a5b17 <= x[5] & y;
	a6b17 <= x[6] & y;
	a7b17 <= x[7] & y;
	a8b17 <= x[8] & y;
	a9b17 <= x[9] & y;
	a10b17 <= x[10] & y;
	a11b17 <= x[11] & y;
	a12b17 <= x[12] & y;
	a13b17 <= x[13] & y;
	a14b17 <= x[14] & y;
	a15b17 <= x[15] & y;
	a16b17 <= x[16] & y;
	a17b17 <= x[17] & y;
	a18b17 <= x[18] & y;
	a19b17 <= x[19] & y;
	a20b17 <= x[20] & y;
	a21b17 <= x[21] & y;
	a22b17 <= x[22] & y;
	a23b17 <= x[23] & y;
	a24b17 <= x[24] & y;
	a25b17 <= x[25] & y;
	a26b17 <= x[26] & y;
	a27b17 <= x[27] & y;
	a28b17 <= x[28] & y;
	a29b17 <= x[29] & y;
	a30b17 <= x[30] & y;
	a31b17 <= x[31] & y;
end

endmodule

module GenPPRow18(x,y,a0b18,a1b18,a2b18,a3b18,a4b18,a5b18,a6b18,a7b18,a8b18,a9b18,a10b18,a11b18,a12b18,a13b18,a14b18,a15b18,a16b18,a17b18,a18b18,a19b18,a20b18,a21b18,a22b18,a23b18,a24b18,a25b18,a26b18,a27b18,a28b18,a29b18,a30b18,a31b18);
input [31:0] x;
input y;
output reg a0b18,a1b18,a2b18,a3b18,a4b18,a5b18,a6b18,a7b18,a8b18,a9b18,a10b18,a11b18,a12b18,a13b18,a14b18,a15b18,a16b18,a17b18,a18b18,a19b18,a20b18,a21b18,a22b18,a23b18,a24b18,a25b18,a26b18,a27b18,a28b18,a29b18,a30b18,a31b18;

always@(x,y)begin
	a0b18 <= x[0] & y;
	a1b18 <= x[1] & y;
	a2b18 <= x[2] & y;
	a3b18 <= x[3] & y;
	a4b18 <= x[4] & y;
	a5b18 <= x[5] & y;
	a6b18 <= x[6] & y;
	a7b18 <= x[7] & y;
	a8b18 <= x[8] & y;
	a9b18 <= x[9] & y;
	a10b18 <= x[10] & y;
	a11b18 <= x[11] & y;
	a12b18 <= x[12] & y;
	a13b18 <= x[13] & y;
	a14b18 <= x[14] & y;
	a15b18 <= x[15] & y;
	a16b18 <= x[16] & y;
	a17b18 <= x[17] & y;
	a18b18 <= x[18] & y;
	a19b18 <= x[19] & y;
	a20b18 <= x[20] & y;
	a21b18 <= x[21] & y;
	a22b18 <= x[22] & y;
	a23b18 <= x[23] & y;
	a24b18 <= x[24] & y;
	a25b18 <= x[25] & y;
	a26b18 <= x[26] & y;
	a27b18 <= x[27] & y;
	a28b18 <= x[28] & y;
	a29b18 <= x[29] & y;
	a30b18 <= x[30] & y;
	a31b18 <= x[31] & y;
end

endmodule

module GenPPRow19(x,y,a0b19,a1b19,a2b19,a3b19,a4b19,a5b19,a6b19,a7b19,a8b19,a9b19,a10b19,a11b19,a12b19,a13b19,a14b19,a15b19,a16b19,a17b19,a18b19,a19b19,a20b19,a21b19,a22b19,a23b19,a24b19,a25b19,a26b19,a27b19,a28b19,a29b19,a30b19,a31b19);
input [31:0] x;
input y;
output reg a0b19,a1b19,a2b19,a3b19,a4b19,a5b19,a6b19,a7b19,a8b19,a9b19,a10b19,a11b19,a12b19,a13b19,a14b19,a15b19,a16b19,a17b19,a18b19,a19b19,a20b19,a21b19,a22b19,a23b19,a24b19,a25b19,a26b19,a27b19,a28b19,a29b19,a30b19,a31b19;

always@(x,y)begin
	a0b19 <= x[0] & y;
	a1b19 <= x[1] & y;
	a2b19 <= x[2] & y;
	a3b19 <= x[3] & y;
	a4b19 <= x[4] & y;
	a5b19 <= x[5] & y;
	a6b19 <= x[6] & y;
	a7b19 <= x[7] & y;
	a8b19 <= x[8] & y;
	a9b19 <= x[9] & y;
	a10b19 <= x[10] & y;
	a11b19 <= x[11] & y;
	a12b19 <= x[12] & y;
	a13b19 <= x[13] & y;
	a14b19 <= x[14] & y;
	a15b19 <= x[15] & y;
	a16b19 <= x[16] & y;
	a17b19 <= x[17] & y;
	a18b19 <= x[18] & y;
	a19b19 <= x[19] & y;
	a20b19 <= x[20] & y;
	a21b19 <= x[21] & y;
	a22b19 <= x[22] & y;
	a23b19 <= x[23] & y;
	a24b19 <= x[24] & y;
	a25b19 <= x[25] & y;
	a26b19 <= x[26] & y;
	a27b19 <= x[27] & y;
	a28b19 <= x[28] & y;
	a29b19 <= x[29] & y;
	a30b19 <= x[30] & y;
	a31b19 <= x[31] & y;
end

endmodule

module GenPPRow20(x,y,a0b20,a1b20,a2b20,a3b20,a4b20,a5b20,a6b20,a7b20,a8b20,a9b20,a10b20,a11b20,a12b20,a13b20,a14b20,a15b20,a16b20,a17b20,a18b20,a19b20,a20b20,a21b20,a22b20,a23b20,a24b20,a25b20,a26b20,a27b20,a28b20,a29b20,a30b20,a31b20);
input [31:0] x;
input y;
output reg a0b20,a1b20,a2b20,a3b20,a4b20,a5b20,a6b20,a7b20,a8b20,a9b20,a10b20,a11b20,a12b20,a13b20,a14b20,a15b20,a16b20,a17b20,a18b20,a19b20,a20b20,a21b20,a22b20,a23b20,a24b20,a25b20,a26b20,a27b20,a28b20,a29b20,a30b20,a31b20;

always@(x,y)begin
	a0b20 <= x[0] & y;
	a1b20 <= x[1] & y;
	a2b20 <= x[2] & y;
	a3b20 <= x[3] & y;
	a4b20 <= x[4] & y;
	a5b20 <= x[5] & y;
	a6b20 <= x[6] & y;
	a7b20 <= x[7] & y;
	a8b20 <= x[8] & y;
	a9b20 <= x[9] & y;
	a10b20 <= x[10] & y;
	a11b20 <= x[11] & y;
	a12b20 <= x[12] & y;
	a13b20 <= x[13] & y;
	a14b20 <= x[14] & y;
	a15b20 <= x[15] & y;
	a16b20 <= x[16] & y;
	a17b20 <= x[17] & y;
	a18b20 <= x[18] & y;
	a19b20 <= x[19] & y;
	a20b20 <= x[20] & y;
	a21b20 <= x[21] & y;
	a22b20 <= x[22] & y;
	a23b20 <= x[23] & y;
	a24b20 <= x[24] & y;
	a25b20 <= x[25] & y;
	a26b20 <= x[26] & y;
	a27b20 <= x[27] & y;
	a28b20 <= x[28] & y;
	a29b20 <= x[29] & y;
	a30b20 <= x[30] & y;
	a31b20 <= x[31] & y;
end

endmodule

module GenPPRow21(x,y,a0b21,a1b21,a2b21,a3b21,a4b21,a5b21,a6b21,a7b21,a8b21,a9b21,a10b21,a11b21,a12b21,a13b21,a14b21,a15b21,a16b21,a17b21,a18b21,a19b21,a20b21,a21b21,a22b21,a23b21,a24b21,a25b21,a26b21,a27b21,a28b21,a29b21,a30b21,a31b21);
input [31:0] x;
input y;
output reg a0b21,a1b21,a2b21,a3b21,a4b21,a5b21,a6b21,a7b21,a8b21,a9b21,a10b21,a11b21,a12b21,a13b21,a14b21,a15b21,a16b21,a17b21,a18b21,a19b21,a20b21,a21b21,a22b21,a23b21,a24b21,a25b21,a26b21,a27b21,a28b21,a29b21,a30b21,a31b21;

always@(x,y)begin
	a0b21 <= x[0] & y;
	a1b21 <= x[1] & y;
	a2b21 <= x[2] & y;
	a3b21 <= x[3] & y;
	a4b21 <= x[4] & y;
	a5b21 <= x[5] & y;
	a6b21 <= x[6] & y;
	a7b21 <= x[7] & y;
	a8b21 <= x[8] & y;
	a9b21 <= x[9] & y;
	a10b21 <= x[10] & y;
	a11b21 <= x[11] & y;
	a12b21 <= x[12] & y;
	a13b21 <= x[13] & y;
	a14b21 <= x[14] & y;
	a15b21 <= x[15] & y;
	a16b21 <= x[16] & y;
	a17b21 <= x[17] & y;
	a18b21 <= x[18] & y;
	a19b21 <= x[19] & y;
	a20b21 <= x[20] & y;
	a21b21 <= x[21] & y;
	a22b21 <= x[22] & y;
	a23b21 <= x[23] & y;
	a24b21 <= x[24] & y;
	a25b21 <= x[25] & y;
	a26b21 <= x[26] & y;
	a27b21 <= x[27] & y;
	a28b21 <= x[28] & y;
	a29b21 <= x[29] & y;
	a30b21 <= x[30] & y;
	a31b21 <= x[31] & y;
end

endmodule

module GenPPRow22(x,y,a0b22,a1b22,a2b22,a3b22,a4b22,a5b22,a6b22,a7b22,a8b22,a9b22,a10b22,a11b22,a12b22,a13b22,a14b22,a15b22,a16b22,a17b22,a18b22,a19b22,a20b22,a21b22,a22b22,a23b22,a24b22,a25b22,a26b22,a27b22,a28b22,a29b22,a30b22,a31b22);
input [31:0] x;
input y;
output reg a0b22,a1b22,a2b22,a3b22,a4b22,a5b22,a6b22,a7b22,a8b22,a9b22,a10b22,a11b22,a12b22,a13b22,a14b22,a15b22,a16b22,a17b22,a18b22,a19b22,a20b22,a21b22,a22b22,a23b22,a24b22,a25b22,a26b22,a27b22,a28b22,a29b22,a30b22,a31b22;

always@(x,y)begin
	a0b22 <= x[0] & y;
	a1b22 <= x[1] & y;
	a2b22 <= x[2] & y;
	a3b22 <= x[3] & y;
	a4b22 <= x[4] & y;
	a5b22 <= x[5] & y;
	a6b22 <= x[6] & y;
	a7b22 <= x[7] & y;
	a8b22 <= x[8] & y;
	a9b22 <= x[9] & y;
	a10b22 <= x[10] & y;
	a11b22 <= x[11] & y;
	a12b22 <= x[12] & y;
	a13b22 <= x[13] & y;
	a14b22 <= x[14] & y;
	a15b22 <= x[15] & y;
	a16b22 <= x[16] & y;
	a17b22 <= x[17] & y;
	a18b22 <= x[18] & y;
	a19b22 <= x[19] & y;
	a20b22 <= x[20] & y;
	a21b22 <= x[21] & y;
	a22b22 <= x[22] & y;
	a23b22 <= x[23] & y;
	a24b22 <= x[24] & y;
	a25b22 <= x[25] & y;
	a26b22 <= x[26] & y;
	a27b22 <= x[27] & y;
	a28b22 <= x[28] & y;
	a29b22 <= x[29] & y;
	a30b22 <= x[30] & y;
	a31b22 <= x[31] & y;
end

endmodule

module GenPPRow23(x,y,a0b23,a1b23,a2b23,a3b23,a4b23,a5b23,a6b23,a7b23,a8b23,a9b23,a10b23,a11b23,a12b23,a13b23,a14b23,a15b23,a16b23,a17b23,a18b23,a19b23,a20b23,a21b23,a22b23,a23b23,a24b23,a25b23,a26b23,a27b23,a28b23,a29b23,a30b23,a31b23);
input [31:0] x;
input y;
output reg a0b23,a1b23,a2b23,a3b23,a4b23,a5b23,a6b23,a7b23,a8b23,a9b23,a10b23,a11b23,a12b23,a13b23,a14b23,a15b23,a16b23,a17b23,a18b23,a19b23,a20b23,a21b23,a22b23,a23b23,a24b23,a25b23,a26b23,a27b23,a28b23,a29b23,a30b23,a31b23;

always@(x,y)begin
	a0b23 <= x[0] & y;
	a1b23 <= x[1] & y;
	a2b23 <= x[2] & y;
	a3b23 <= x[3] & y;
	a4b23 <= x[4] & y;
	a5b23 <= x[5] & y;
	a6b23 <= x[6] & y;
	a7b23 <= x[7] & y;
	a8b23 <= x[8] & y;
	a9b23 <= x[9] & y;
	a10b23 <= x[10] & y;
	a11b23 <= x[11] & y;
	a12b23 <= x[12] & y;
	a13b23 <= x[13] & y;
	a14b23 <= x[14] & y;
	a15b23 <= x[15] & y;
	a16b23 <= x[16] & y;
	a17b23 <= x[17] & y;
	a18b23 <= x[18] & y;
	a19b23 <= x[19] & y;
	a20b23 <= x[20] & y;
	a21b23 <= x[21] & y;
	a22b23 <= x[22] & y;
	a23b23 <= x[23] & y;
	a24b23 <= x[24] & y;
	a25b23 <= x[25] & y;
	a26b23 <= x[26] & y;
	a27b23 <= x[27] & y;
	a28b23 <= x[28] & y;
	a29b23 <= x[29] & y;
	a30b23 <= x[30] & y;
	a31b23 <= x[31] & y;
end

endmodule

module GenPPRow24(x,y,a0b24,a1b24,a2b24,a3b24,a4b24,a5b24,a6b24,a7b24,a8b24,a9b24,a10b24,a11b24,a12b24,a13b24,a14b24,a15b24,a16b24,a17b24,a18b24,a19b24,a20b24,a21b24,a22b24,a23b24,a24b24,a25b24,a26b24,a27b24,a28b24,a29b24,a30b24,a31b24);
input [31:0] x;
input y;
output reg a0b24,a1b24,a2b24,a3b24,a4b24,a5b24,a6b24,a7b24,a8b24,a9b24,a10b24,a11b24,a12b24,a13b24,a14b24,a15b24,a16b24,a17b24,a18b24,a19b24,a20b24,a21b24,a22b24,a23b24,a24b24,a25b24,a26b24,a27b24,a28b24,a29b24,a30b24,a31b24;

always@(x,y)begin
	a0b24 <= x[0] & y;
	a1b24 <= x[1] & y;
	a2b24 <= x[2] & y;
	a3b24 <= x[3] & y;
	a4b24 <= x[4] & y;
	a5b24 <= x[5] & y;
	a6b24 <= x[6] & y;
	a7b24 <= x[7] & y;
	a8b24 <= x[8] & y;
	a9b24 <= x[9] & y;
	a10b24 <= x[10] & y;
	a11b24 <= x[11] & y;
	a12b24 <= x[12] & y;
	a13b24 <= x[13] & y;
	a14b24 <= x[14] & y;
	a15b24 <= x[15] & y;
	a16b24 <= x[16] & y;
	a17b24 <= x[17] & y;
	a18b24 <= x[18] & y;
	a19b24 <= x[19] & y;
	a20b24 <= x[20] & y;
	a21b24 <= x[21] & y;
	a22b24 <= x[22] & y;
	a23b24 <= x[23] & y;
	a24b24 <= x[24] & y;
	a25b24 <= x[25] & y;
	a26b24 <= x[26] & y;
	a27b24 <= x[27] & y;
	a28b24 <= x[28] & y;
	a29b24 <= x[29] & y;
	a30b24 <= x[30] & y;
	a31b24 <= x[31] & y;
end

endmodule

module GenPPRow25(x,y,a0b25,a1b25,a2b25,a3b25,a4b25,a5b25,a6b25,a7b25,a8b25,a9b25,a10b25,a11b25,a12b25,a13b25,a14b25,a15b25,a16b25,a17b25,a18b25,a19b25,a20b25,a21b25,a22b25,a23b25,a24b25,a25b25,a26b25,a27b25,a28b25,a29b25,a30b25,a31b25);
input [31:0] x;
input y;
output reg a0b25,a1b25,a2b25,a3b25,a4b25,a5b25,a6b25,a7b25,a8b25,a9b25,a10b25,a11b25,a12b25,a13b25,a14b25,a15b25,a16b25,a17b25,a18b25,a19b25,a20b25,a21b25,a22b25,a23b25,a24b25,a25b25,a26b25,a27b25,a28b25,a29b25,a30b25,a31b25;

always@(x,y)begin
	a0b25 <= x[0] & y;
	a1b25 <= x[1] & y;
	a2b25 <= x[2] & y;
	a3b25 <= x[3] & y;
	a4b25 <= x[4] & y;
	a5b25 <= x[5] & y;
	a6b25 <= x[6] & y;
	a7b25 <= x[7] & y;
	a8b25 <= x[8] & y;
	a9b25 <= x[9] & y;
	a10b25 <= x[10] & y;
	a11b25 <= x[11] & y;
	a12b25 <= x[12] & y;
	a13b25 <= x[13] & y;
	a14b25 <= x[14] & y;
	a15b25 <= x[15] & y;
	a16b25 <= x[16] & y;
	a17b25 <= x[17] & y;
	a18b25 <= x[18] & y;
	a19b25 <= x[19] & y;
	a20b25 <= x[20] & y;
	a21b25 <= x[21] & y;
	a22b25 <= x[22] & y;
	a23b25 <= x[23] & y;
	a24b25 <= x[24] & y;
	a25b25 <= x[25] & y;
	a26b25 <= x[26] & y;
	a27b25 <= x[27] & y;
	a28b25 <= x[28] & y;
	a29b25 <= x[29] & y;
	a30b25 <= x[30] & y;
	a31b25 <= x[31] & y;
end

endmodule

module GenPPRow26(x,y,a0b26,a1b26,a2b26,a3b26,a4b26,a5b26,a6b26,a7b26,a8b26,a9b26,a10b26,a11b26,a12b26,a13b26,a14b26,a15b26,a16b26,a17b26,a18b26,a19b26,a20b26,a21b26,a22b26,a23b26,a24b26,a25b26,a26b26,a27b26,a28b26,a29b26,a30b26,a31b26);
input [31:0] x;
input y;
output reg a0b26,a1b26,a2b26,a3b26,a4b26,a5b26,a6b26,a7b26,a8b26,a9b26,a10b26,a11b26,a12b26,a13b26,a14b26,a15b26,a16b26,a17b26,a18b26,a19b26,a20b26,a21b26,a22b26,a23b26,a24b26,a25b26,a26b26,a27b26,a28b26,a29b26,a30b26,a31b26;

always@(x,y)begin
	a0b26 <= x[0] & y;
	a1b26 <= x[1] & y;
	a2b26 <= x[2] & y;
	a3b26 <= x[3] & y;
	a4b26 <= x[4] & y;
	a5b26 <= x[5] & y;
	a6b26 <= x[6] & y;
	a7b26 <= x[7] & y;
	a8b26 <= x[8] & y;
	a9b26 <= x[9] & y;
	a10b26 <= x[10] & y;
	a11b26 <= x[11] & y;
	a12b26 <= x[12] & y;
	a13b26 <= x[13] & y;
	a14b26 <= x[14] & y;
	a15b26 <= x[15] & y;
	a16b26 <= x[16] & y;
	a17b26 <= x[17] & y;
	a18b26 <= x[18] & y;
	a19b26 <= x[19] & y;
	a20b26 <= x[20] & y;
	a21b26 <= x[21] & y;
	a22b26 <= x[22] & y;
	a23b26 <= x[23] & y;
	a24b26 <= x[24] & y;
	a25b26 <= x[25] & y;
	a26b26 <= x[26] & y;
	a27b26 <= x[27] & y;
	a28b26 <= x[28] & y;
	a29b26 <= x[29] & y;
	a30b26 <= x[30] & y;
	a31b26 <= x[31] & y;
end

endmodule

module GenPPRow27(x,y,a0b27,a1b27,a2b27,a3b27,a4b27,a5b27,a6b27,a7b27,a8b27,a9b27,a10b27,a11b27,a12b27,a13b27,a14b27,a15b27,a16b27,a17b27,a18b27,a19b27,a20b27,a21b27,a22b27,a23b27,a24b27,a25b27,a26b27,a27b27,a28b27,a29b27,a30b27,a31b27);
input [31:0] x;
input y;
output reg a0b27,a1b27,a2b27,a3b27,a4b27,a5b27,a6b27,a7b27,a8b27,a9b27,a10b27,a11b27,a12b27,a13b27,a14b27,a15b27,a16b27,a17b27,a18b27,a19b27,a20b27,a21b27,a22b27,a23b27,a24b27,a25b27,a26b27,a27b27,a28b27,a29b27,a30b27,a31b27;

always@(x,y)begin
	a0b27 <= x[0] & y;
	a1b27 <= x[1] & y;
	a2b27 <= x[2] & y;
	a3b27 <= x[3] & y;
	a4b27 <= x[4] & y;
	a5b27 <= x[5] & y;
	a6b27 <= x[6] & y;
	a7b27 <= x[7] & y;
	a8b27 <= x[8] & y;
	a9b27 <= x[9] & y;
	a10b27 <= x[10] & y;
	a11b27 <= x[11] & y;
	a12b27 <= x[12] & y;
	a13b27 <= x[13] & y;
	a14b27 <= x[14] & y;
	a15b27 <= x[15] & y;
	a16b27 <= x[16] & y;
	a17b27 <= x[17] & y;
	a18b27 <= x[18] & y;
	a19b27 <= x[19] & y;
	a20b27 <= x[20] & y;
	a21b27 <= x[21] & y;
	a22b27 <= x[22] & y;
	a23b27 <= x[23] & y;
	a24b27 <= x[24] & y;
	a25b27 <= x[25] & y;
	a26b27 <= x[26] & y;
	a27b27 <= x[27] & y;
	a28b27 <= x[28] & y;
	a29b27 <= x[29] & y;
	a30b27 <= x[30] & y;
	a31b27 <= x[31] & y;
end

endmodule

module GenPPRow28(x,y,a0b28,a1b28,a2b28,a3b28,a4b28,a5b28,a6b28,a7b28,a8b28,a9b28,a10b28,a11b28,a12b28,a13b28,a14b28,a15b28,a16b28,a17b28,a18b28,a19b28,a20b28,a21b28,a22b28,a23b28,a24b28,a25b28,a26b28,a27b28,a28b28,a29b28,a30b28,a31b28);
input [31:0] x;
input y;
output reg a0b28,a1b28,a2b28,a3b28,a4b28,a5b28,a6b28,a7b28,a8b28,a9b28,a10b28,a11b28,a12b28,a13b28,a14b28,a15b28,a16b28,a17b28,a18b28,a19b28,a20b28,a21b28,a22b28,a23b28,a24b28,a25b28,a26b28,a27b28,a28b28,a29b28,a30b28,a31b28;

always@(x,y)begin
	a0b28 <= x[0] & y;
	a1b28 <= x[1] & y;
	a2b28 <= x[2] & y;
	a3b28 <= x[3] & y;
	a4b28 <= x[4] & y;
	a5b28 <= x[5] & y;
	a6b28 <= x[6] & y;
	a7b28 <= x[7] & y;
	a8b28 <= x[8] & y;
	a9b28 <= x[9] & y;
	a10b28 <= x[10] & y;
	a11b28 <= x[11] & y;
	a12b28 <= x[12] & y;
	a13b28 <= x[13] & y;
	a14b28 <= x[14] & y;
	a15b28 <= x[15] & y;
	a16b28 <= x[16] & y;
	a17b28 <= x[17] & y;
	a18b28 <= x[18] & y;
	a19b28 <= x[19] & y;
	a20b28 <= x[20] & y;
	a21b28 <= x[21] & y;
	a22b28 <= x[22] & y;
	a23b28 <= x[23] & y;
	a24b28 <= x[24] & y;
	a25b28 <= x[25] & y;
	a26b28 <= x[26] & y;
	a27b28 <= x[27] & y;
	a28b28 <= x[28] & y;
	a29b28 <= x[29] & y;
	a30b28 <= x[30] & y;
	a31b28 <= x[31] & y;
end

endmodule

module GenPPRow29(x,y,a0b29,a1b29,a2b29,a3b29,a4b29,a5b29,a6b29,a7b29,a8b29,a9b29,a10b29,a11b29,a12b29,a13b29,a14b29,a15b29,a16b29,a17b29,a18b29,a19b29,a20b29,a21b29,a22b29,a23b29,a24b29,a25b29,a26b29,a27b29,a28b29,a29b29,a30b29,a31b29);
input [31:0] x;
input y;
output reg a0b29,a1b29,a2b29,a3b29,a4b29,a5b29,a6b29,a7b29,a8b29,a9b29,a10b29,a11b29,a12b29,a13b29,a14b29,a15b29,a16b29,a17b29,a18b29,a19b29,a20b29,a21b29,a22b29,a23b29,a24b29,a25b29,a26b29,a27b29,a28b29,a29b29,a30b29,a31b29;

always@(x,y)begin
	a0b29 <= x[0] & y;
	a1b29 <= x[1] & y;
	a2b29 <= x[2] & y;
	a3b29 <= x[3] & y;
	a4b29 <= x[4] & y;
	a5b29 <= x[5] & y;
	a6b29 <= x[6] & y;
	a7b29 <= x[7] & y;
	a8b29 <= x[8] & y;
	a9b29 <= x[9] & y;
	a10b29 <= x[10] & y;
	a11b29 <= x[11] & y;
	a12b29 <= x[12] & y;
	a13b29 <= x[13] & y;
	a14b29 <= x[14] & y;
	a15b29 <= x[15] & y;
	a16b29 <= x[16] & y;
	a17b29 <= x[17] & y;
	a18b29 <= x[18] & y;
	a19b29 <= x[19] & y;
	a20b29 <= x[20] & y;
	a21b29 <= x[21] & y;
	a22b29 <= x[22] & y;
	a23b29 <= x[23] & y;
	a24b29 <= x[24] & y;
	a25b29 <= x[25] & y;
	a26b29 <= x[26] & y;
	a27b29 <= x[27] & y;
	a28b29 <= x[28] & y;
	a29b29 <= x[29] & y;
	a30b29 <= x[30] & y;
	a31b29 <= x[31] & y;
end

endmodule

module GenPPRow30(x,y,a0b30,a1b30,a2b30,a3b30,a4b30,a5b30,a6b30,a7b30,a8b30,a9b30,a10b30,a11b30,a12b30,a13b30,a14b30,a15b30,a16b30,a17b30,a18b30,a19b30,a20b30,a21b30,a22b30,a23b30,a24b30,a25b30,a26b30,a27b30,a28b30,a29b30,a30b30,a31b30);
input [31:0] x;
input y;
output reg a0b30,a1b30,a2b30,a3b30,a4b30,a5b30,a6b30,a7b30,a8b30,a9b30,a10b30,a11b30,a12b30,a13b30,a14b30,a15b30,a16b30,a17b30,a18b30,a19b30,a20b30,a21b30,a22b30,a23b30,a24b30,a25b30,a26b30,a27b30,a28b30,a29b30,a30b30,a31b30;

always@(x,y)begin
	a0b30 <= x[0] & y;
	a1b30 <= x[1] & y;
	a2b30 <= x[2] & y;
	a3b30 <= x[3] & y;
	a4b30 <= x[4] & y;
	a5b30 <= x[5] & y;
	a6b30 <= x[6] & y;
	a7b30 <= x[7] & y;
	a8b30 <= x[8] & y;
	a9b30 <= x[9] & y;
	a10b30 <= x[10] & y;
	a11b30 <= x[11] & y;
	a12b30 <= x[12] & y;
	a13b30 <= x[13] & y;
	a14b30 <= x[14] & y;
	a15b30 <= x[15] & y;
	a16b30 <= x[16] & y;
	a17b30 <= x[17] & y;
	a18b30 <= x[18] & y;
	a19b30 <= x[19] & y;
	a20b30 <= x[20] & y;
	a21b30 <= x[21] & y;
	a22b30 <= x[22] & y;
	a23b30 <= x[23] & y;
	a24b30 <= x[24] & y;
	a25b30 <= x[25] & y;
	a26b30 <= x[26] & y;
	a27b30 <= x[27] & y;
	a28b30 <= x[28] & y;
	a29b30 <= x[29] & y;
	a30b30 <= x[30] & y;
	a31b30 <= x[31] & y;
end

endmodule

module GenPPRow31(x,y,a0b31,a1b31,a2b31,a3b31,a4b31,a5b31,a6b31,a7b31,a8b31,a9b31,a10b31,a11b31,a12b31,a13b31,a14b31,a15b31,a16b31,a17b31,a18b31,a19b31,a20b31,a21b31,a22b31,a23b31,a24b31,a25b31,a26b31,a27b31,a28b31,a29b31,a30b31,a31b31);
input [31:0] x;
input y;
output reg a0b31,a1b31,a2b31,a3b31,a4b31,a5b31,a6b31,a7b31,a8b31,a9b31,a10b31,a11b31,a12b31,a13b31,a14b31,a15b31,a16b31,a17b31,a18b31,a19b31,a20b31,a21b31,a22b31,a23b31,a24b31,a25b31,a26b31,a27b31,a28b31,a29b31,a30b31,a31b31;

always@(x,y)begin
	a0b31 <= x[0] & y;
	a1b31 <= x[1] & y;
	a2b31 <= x[2] & y;
	a3b31 <= x[3] & y;
	a4b31 <= x[4] & y;
	a5b31 <= x[5] & y;
	a6b31 <= x[6] & y;
	a7b31 <= x[7] & y;
	a8b31 <= x[8] & y;
	a9b31 <= x[9] & y;
	a10b31 <= x[10] & y;
	a11b31 <= x[11] & y;
	a12b31 <= x[12] & y;
	a13b31 <= x[13] & y;
	a14b31 <= x[14] & y;
	a15b31 <= x[15] & y;
	a16b31 <= x[16] & y;
	a17b31 <= x[17] & y;
	a18b31 <= x[18] & y;
	a19b31 <= x[19] & y;
	a20b31 <= x[20] & y;
	a21b31 <= x[21] & y;
	a22b31 <= x[22] & y;
	a23b31 <= x[23] & y;
	a24b31 <= x[24] & y;
	a25b31 <= x[25] & y;
	a26b31 <= x[26] & y;
	a27b31 <= x[27] & y;
	a28b31 <= x[28] & y;
	a29b31 <= x[29] & y;
	a30b31 <= x[30] & y;
	a31b31 <= x[31] & y;
end

endmodule
