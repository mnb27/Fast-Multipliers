`timescale 1ns / 1ps

module stage0(r0,r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16,r17,r18,r19,r20,r21,r22,r23,r24,r25,r26,r27,r28,r29,r30,r31,r32,r33,r34,r35,r36,r37,r38,r39,r40,r41,r42,r43,r44,r45,r46,r47,r48,r49,r50,r51,r52,r53,r54,r55,r56,r57,r58,r59,r60,r61,r62,r63,r64,r65,r66,r67,r68,r69,r70,r71,r72,r73,r74,r75,r76,r77,r78,r79,r80,r81,r82,r83,r84,r85,r86,r87,r88,r89,r90,r91,r92,r93,r94,r95,r96,r97,r98,r99,r100,r101,r102,r103,r104,r105,r106,r107,r108,r109,r110,r111,r112,r113,r114,r115,r116,r117,r118,r119,r120,r121,r122,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,s61,p2,p64);
input r0,r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16,r17,r18,r19,r20,r21,r22,r23,r24,r25,r26,r27,r28,r29,r30,r31,r32,r33,r34,r35,r36,r37,r38,r39,r40,r41,r42,r43,r44,r45,r46,r47,r48,r49,r50,r51,r52,r53,r54,r55,r56,r57,r58,r59,r60,r61,r62,r63,r64,r65,r66,r67,r68,r69,r70,r71,r72,r73,r74,r75,r76,r77,r78,r79,r80,r81,r82,r83,r84,r85,r86,r87,r88,r89,r90,r91,r92,r93,r94,r95,r96,r97,r98,r99,r100,r101,r102,r103,r104,r105,r106,r107,r108,r109,r110,r111,r112,r113,r114,r115,r116,r117,r118,r119,r120,r121,r122;
output s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,s61,p2,p64;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,d49,d50,d51,d52,d53,d54,d55,d56,d57,d58,d59,d60,d61;


full_adder fa0(r0,r62,1'b0,p2,d1);
full_adder fa1(r1,r63,d1,s1,d2);
full_adder fa2(r2,r64,d2,s2,d3);
full_adder fa3(r3,r65,d3,s3,d4);
full_adder fa4(r4,r66,d4,s4,d5);
full_adder fa5(r5,r67,d5,s5,d6);
full_adder fa6(r6,r68,d6,s6,d7);
full_adder fa7(r7,r69,d7,s7,d8);
full_adder fa8(r8,r70,d8,s8,d9);
full_adder fa9(r9,r71,d9,s9,d10);
full_adder fa10(r10,r72,d10,s10,d11);
full_adder fa11(r11,r73,d11,s11,d12);
full_adder fa12(r12,r74,d12,s12,d13);
full_adder fa13(r13,r75,d13,s13,d14);
full_adder fa14(r14,r76,d14,s14,d15);
full_adder fa15(r15,r77,d15,s15,d16);
full_adder fa16(r16,r78,d16,s16,d17);
full_adder fa17(r17,r79,d17,s17,d18);
full_adder fa18(r18,r80,d18,s18,d19);
full_adder fa19(r19,r81,d19,s19,d20);
full_adder fa20(r20,r82,d20,s20,d21);
full_adder fa21(r21,r83,d21,s21,d22);
full_adder fa22(r22,r84,d22,s22,d23);
full_adder fa23(r23,r85,d23,s23,d24);
full_adder fa24(r24,r86,d24,s24,d25);
full_adder fa25(r25,r87,d25,s25,d26);
full_adder fa26(r26,r88,d26,s26,d27);
full_adder fa27(r27,r89,d27,s27,d28);
full_adder fa28(r28,r90,d28,s28,d29);
full_adder fa29(r29,r91,d29,s29,d30);
full_adder fa30(r30,r92,d30,s30,d31);
full_adder fa31(r31,r93,d31,s31,d32);
full_adder fa32(r32,r94,d32,s32,d33);
full_adder fa33(r33,r95,d33,s33,d34);
full_adder fa34(r34,r96,d34,s34,d35);
full_adder fa35(r35,r97,d35,s35,d36);
full_adder fa36(r36,r98,d36,s36,d37);
full_adder fa37(r37,r99,d37,s37,d38);
full_adder fa38(r38,r100,d38,s38,d39);
full_adder fa39(r39,r101,d39,s39,d40);
full_adder fa40(r40,r102,d40,s40,d41);
full_adder fa41(r41,r103,d41,s41,d42);
full_adder fa42(r42,r104,d42,s42,d43);
full_adder fa43(r43,r105,d43,s43,d44);
full_adder fa44(r44,r106,d44,s44,d45);
full_adder fa45(r45,r107,d45,s45,d46);
full_adder fa46(r46,r108,d46,s46,d47);
full_adder fa47(r47,r109,d47,s47,d48);
full_adder fa48(r48,r110,d48,s48,d49);
full_adder fa49(r49,r111,d49,s49,d50);
full_adder fa50(r50,r112,d50,s50,d51);
full_adder fa51(r51,r113,d51,s51,d52);
full_adder fa52(r52,r114,d52,s52,d53);
full_adder fa53(r53,r115,d53,s53,d54);
full_adder fa54(r54,r116,d54,s54,d55);
full_adder fa55(r55,r117,d55,s55,d56);
full_adder fa56(r56,r118,d56,s56,d57);
full_adder fa57(r57,r119,d57,s57,d58);
full_adder fa58(r58,r120,d58,s58,d59);
full_adder fa59(r59,r121,d59,s59,d60);
full_adder fa60(r60,r122,d60,s60,d61);
full_adder fa61(r61,1'b0,d61,s61,p64);

endmodule

module stage1(r123,r124,r125,r126,r127,r128,r129,r130,r131,r132,r133,r134,r135,r136,r137,r138,r139,r140,r141,r142,r143,r144,r145,r146,r147,r148,r149,r150,r151,r152,r153,r154,r155,r156,r157,r158,r159,r160,r161,r162,r163,r164,r165,r166,r167,r168,r169,r170,r171,r172,r173,r174,r175,r176,r177,r178,r179,r180,r181,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,s61,s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74,s75,s76,s77,s78,s79,s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s90,s91,s92,s93,s94,s95,s96,s97,s98,s99,s100,s101,s102,s103,s104,s105,s106,s107,s108,s109,s110,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120,p3,p63);
input r123,r124,r125,r126,r127,r128,r129,r130,r131,r132,r133,r134,r135,r136,r137,r138,r139,r140,r141,r142,r143,r144,r145,r146,r147,r148,r149,r150,r151,r152,r153,r154,r155,r156,r157,r158,r159,r160,r161,r162,r163,r164,r165,r166,r167,r168,r169,r170,r171,r172,r173,r174,r175,r176,r177,r178,r179,r180,r181,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,s61;
output s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74,s75,s76,s77,s78,s79,s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s90,s91,s92,s93,s94,s95,s96,s97,s98,s99,s100,s101,s102,s103,s104,s105,s106,s107,s108,s109,s110,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120,p3,p63;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,d49,d50,d51,d52,d53,d54,d55,d56,d57,d58,d59,d60;


full_adder fa0(s1,r123,1'b0,p3,d1);
full_adder fa1(s2,r124,d1,s62,d2);
full_adder fa2(s3,r125,d2,s63,d3);
full_adder fa3(s4,r126,d3,s64,d4);
full_adder fa4(s5,r127,d4,s65,d5);
full_adder fa5(s6,r128,d5,s66,d6);
full_adder fa6(s7,r129,d6,s67,d7);
full_adder fa7(s8,r130,d7,s68,d8);
full_adder fa8(s9,r131,d8,s69,d9);
full_adder fa9(s10,r132,d9,s70,d10);
full_adder fa10(s11,r133,d10,s71,d11);
full_adder fa11(s12,r134,d11,s72,d12);
full_adder fa12(s13,r135,d12,s73,d13);
full_adder fa13(s14,r136,d13,s74,d14);
full_adder fa14(s15,r137,d14,s75,d15);
full_adder fa15(s16,r138,d15,s76,d16);
full_adder fa16(s17,r139,d16,s77,d17);
full_adder fa17(s18,r140,d17,s78,d18);
full_adder fa18(s19,r141,d18,s79,d19);
full_adder fa19(s20,r142,d19,s80,d20);
full_adder fa20(s21,r143,d20,s81,d21);
full_adder fa21(s22,r144,d21,s82,d22);
full_adder fa22(s23,r145,d22,s83,d23);
full_adder fa23(s24,r146,d23,s84,d24);
full_adder fa24(s25,r147,d24,s85,d25);
full_adder fa25(s26,r148,d25,s86,d26);
full_adder fa26(s27,r149,d26,s87,d27);
full_adder fa27(s28,r150,d27,s88,d28);
full_adder fa28(s29,r151,d28,s89,d29);
full_adder fa29(s30,r152,d29,s90,d30);
full_adder fa30(s31,r153,d30,s91,d31);
full_adder fa31(s32,r154,d31,s92,d32);
full_adder fa32(s33,r155,d32,s93,d33);
full_adder fa33(s34,r156,d33,s94,d34);
full_adder fa34(s35,r157,d34,s95,d35);
full_adder fa35(s36,r158,d35,s96,d36);
full_adder fa36(s37,r159,d36,s97,d37);
full_adder fa37(s38,r160,d37,s98,d38);
full_adder fa38(s39,r161,d38,s99,d39);
full_adder fa39(s40,r162,d39,s100,d40);
full_adder fa40(s41,r163,d40,s101,d41);
full_adder fa41(s42,r164,d41,s102,d42);
full_adder fa42(s43,r165,d42,s103,d43);
full_adder fa43(s44,r166,d43,s104,d44);
full_adder fa44(s45,r167,d44,s105,d45);
full_adder fa45(s46,r168,d45,s106,d46);
full_adder fa46(s47,r169,d46,s107,d47);
full_adder fa47(s48,r170,d47,s108,d48);
full_adder fa48(s49,r171,d48,s109,d49);
full_adder fa49(s50,r172,d49,s110,d50);
full_adder fa50(s51,r173,d50,s111,d51);
full_adder fa51(s52,r174,d51,s112,d52);
full_adder fa52(s53,r175,d52,s113,d53);
full_adder fa53(s54,r176,d53,s114,d54);
full_adder fa54(s55,r177,d54,s115,d55);
full_adder fa55(s56,r178,d55,s116,d56);
full_adder fa56(s57,r179,d56,s117,d57);
full_adder fa57(s58,r180,d57,s118,d58);
full_adder fa58(s59,r181,d58,s119,d59);
full_adder fa59(s60,1'b0,d59,s120,d60);
full_adder fa60(s61,1'b0,d60,p63,);

endmodule

module stage2(r182,r183,r184,r185,r186,r187,r188,r189,r190,r191,r192,r193,r194,r195,r196,r197,r198,r199,r200,r201,r202,r203,r204,r205,r206,r207,r208,r209,r210,r211,r212,r213,r214,r215,r216,r217,r218,r219,r220,r221,r222,r223,r224,r225,r226,r227,r228,r229,r230,r231,r232,r233,r234,r235,r236,r237,r238,s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74,s75,s76,s77,s78,s79,s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s90,s91,s92,s93,s94,s95,s96,s97,s98,s99,s100,s101,s102,s103,s104,s105,s106,s107,s108,s109,s110,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120,s121,s122,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s133,s134,s135,s136,s137,s138,s139,s140,s141,s142,s143,s144,s145,s146,s147,s148,s149,s150,s151,s152,s153,s154,s155,s156,s157,s158,s159,s160,s161,s162,s163,s164,s165,s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177,p4,p62);
input r182,r183,r184,r185,r186,r187,r188,r189,r190,r191,r192,r193,r194,r195,r196,r197,r198,r199,r200,r201,r202,r203,r204,r205,r206,r207,r208,r209,r210,r211,r212,r213,r214,r215,r216,r217,r218,r219,r220,r221,r222,r223,r224,r225,r226,r227,r228,r229,r230,r231,r232,r233,r234,r235,r236,r237,r238,s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74,s75,s76,s77,s78,s79,s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s90,s91,s92,s93,s94,s95,s96,s97,s98,s99,s100,s101,s102,s103,s104,s105,s106,s107,s108,s109,s110,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120;
output s121,s122,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s133,s134,s135,s136,s137,s138,s139,s140,s141,s142,s143,s144,s145,s146,s147,s148,s149,s150,s151,s152,s153,s154,s155,s156,s157,s158,s159,s160,s161,s162,s163,s164,s165,s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177,p4,p62;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,d49,d50,d51,d52,d53,d54,d55,d56,d57,d58;


full_adder fa0(s62,r182,1'b0,p4,d1);
full_adder fa1(s63,r183,d1,s121,d2);
full_adder fa2(s64,r184,d2,s122,d3);
full_adder fa3(s65,r185,d3,s123,d4);
full_adder fa4(s66,r186,d4,s124,d5);
full_adder fa5(s67,r187,d5,s125,d6);
full_adder fa6(s68,r188,d6,s126,d7);
full_adder fa7(s69,r189,d7,s127,d8);
full_adder fa8(s70,r190,d8,s128,d9);
full_adder fa9(s71,r191,d9,s129,d10);
full_adder fa10(s72,r192,d10,s130,d11);
full_adder fa11(s73,r193,d11,s131,d12);
full_adder fa12(s74,r194,d12,s132,d13);
full_adder fa13(s75,r195,d13,s133,d14);
full_adder fa14(s76,r196,d14,s134,d15);
full_adder fa15(s77,r197,d15,s135,d16);
full_adder fa16(s78,r198,d16,s136,d17);
full_adder fa17(s79,r199,d17,s137,d18);
full_adder fa18(s80,r200,d18,s138,d19);
full_adder fa19(s81,r201,d19,s139,d20);
full_adder fa20(s82,r202,d20,s140,d21);
full_adder fa21(s83,r203,d21,s141,d22);
full_adder fa22(s84,r204,d22,s142,d23);
full_adder fa23(s85,r205,d23,s143,d24);
full_adder fa24(s86,r206,d24,s144,d25);
full_adder fa25(s87,r207,d25,s145,d26);
full_adder fa26(s88,r208,d26,s146,d27);
full_adder fa27(s89,r209,d27,s147,d28);
full_adder fa28(s90,r210,d28,s148,d29);
full_adder fa29(s91,r211,d29,s149,d30);
full_adder fa30(s92,r212,d30,s150,d31);
full_adder fa31(s93,r213,d31,s151,d32);
full_adder fa32(s94,r214,d32,s152,d33);
full_adder fa33(s95,r215,d33,s153,d34);
full_adder fa34(s96,r216,d34,s154,d35);
full_adder fa35(s97,r217,d35,s155,d36);
full_adder fa36(s98,r218,d36,s156,d37);
full_adder fa37(s99,r219,d37,s157,d38);
full_adder fa38(s100,r220,d38,s158,d39);
full_adder fa39(s101,r221,d39,s159,d40);
full_adder fa40(s102,r222,d40,s160,d41);
full_adder fa41(s103,r223,d41,s161,d42);
full_adder fa42(s104,r224,d42,s162,d43);
full_adder fa43(s105,r225,d43,s163,d44);
full_adder fa44(s106,r226,d44,s164,d45);
full_adder fa45(s107,r227,d45,s165,d46);
full_adder fa46(s108,r228,d46,s166,d47);
full_adder fa47(s109,r229,d47,s167,d48);
full_adder fa48(s110,r230,d48,s168,d49);
full_adder fa49(s111,r231,d49,s169,d50);
full_adder fa50(s112,r232,d50,s170,d51);
full_adder fa51(s113,r233,d51,s171,d52);
full_adder fa52(s114,r234,d52,s172,d53);
full_adder fa53(s115,r235,d53,s173,d54);
full_adder fa54(s116,r236,d54,s174,d55);
full_adder fa55(s117,r237,d55,s175,d56);
full_adder fa56(s118,r238,d56,s176,d57);
full_adder fa57(s119,1'b0,d57,s177,d58);
full_adder fa58(s120,1'b0,d58,p62,);

endmodule

module stage3(r239,r240,r241,r242,r243,r244,r245,r246,r247,r248,r249,r250,r251,r252,r253,r254,r255,r256,r257,r258,r259,r260,r261,r262,r263,r264,r265,r266,r267,r268,r269,r270,r271,r272,r273,r274,r275,r276,r277,r278,r279,r280,r281,r282,r283,r284,r285,r286,r287,r288,r289,r290,r291,r292,r293,s121,s122,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s133,s134,s135,s136,s137,s138,s139,s140,s141,s142,s143,s144,s145,s146,s147,s148,s149,s150,s151,s152,s153,s154,s155,s156,s157,s158,s159,s160,s161,s162,s163,s164,s165,s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177,s178,s179,s180,s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,s226,s227,s228,s229,s230,s231,s232,p5,p61);
input r239,r240,r241,r242,r243,r244,r245,r246,r247,r248,r249,r250,r251,r252,r253,r254,r255,r256,r257,r258,r259,r260,r261,r262,r263,r264,r265,r266,r267,r268,r269,r270,r271,r272,r273,r274,r275,r276,r277,r278,r279,r280,r281,r282,r283,r284,r285,r286,r287,r288,r289,r290,r291,r292,r293,s121,s122,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s133,s134,s135,s136,s137,s138,s139,s140,s141,s142,s143,s144,s145,s146,s147,s148,s149,s150,s151,s152,s153,s154,s155,s156,s157,s158,s159,s160,s161,s162,s163,s164,s165,s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177;
output s178,s179,s180,s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,s226,s227,s228,s229,s230,s231,s232,p5,p61;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,d49,d50,d51,d52,d53,d54,d55,d56;


full_adder fa0(s121,r239,1'b0,p5,d1);
full_adder fa1(s122,r240,d1,s178,d2);
full_adder fa2(s123,r241,d2,s179,d3);
full_adder fa3(s124,r242,d3,s180,d4);
full_adder fa4(s125,r243,d4,s181,d5);
full_adder fa5(s126,r244,d5,s182,d6);
full_adder fa6(s127,r245,d6,s183,d7);
full_adder fa7(s128,r246,d7,s184,d8);
full_adder fa8(s129,r247,d8,s185,d9);
full_adder fa9(s130,r248,d9,s186,d10);
full_adder fa10(s131,r249,d10,s187,d11);
full_adder fa11(s132,r250,d11,s188,d12);
full_adder fa12(s133,r251,d12,s189,d13);
full_adder fa13(s134,r252,d13,s190,d14);
full_adder fa14(s135,r253,d14,s191,d15);
full_adder fa15(s136,r254,d15,s192,d16);
full_adder fa16(s137,r255,d16,s193,d17);
full_adder fa17(s138,r256,d17,s194,d18);
full_adder fa18(s139,r257,d18,s195,d19);
full_adder fa19(s140,r258,d19,s196,d20);
full_adder fa20(s141,r259,d20,s197,d21);
full_adder fa21(s142,r260,d21,s198,d22);
full_adder fa22(s143,r261,d22,s199,d23);
full_adder fa23(s144,r262,d23,s200,d24);
full_adder fa24(s145,r263,d24,s201,d25);
full_adder fa25(s146,r264,d25,s202,d26);
full_adder fa26(s147,r265,d26,s203,d27);
full_adder fa27(s148,r266,d27,s204,d28);
full_adder fa28(s149,r267,d28,s205,d29);
full_adder fa29(s150,r268,d29,s206,d30);
full_adder fa30(s151,r269,d30,s207,d31);
full_adder fa31(s152,r270,d31,s208,d32);
full_adder fa32(s153,r271,d32,s209,d33);
full_adder fa33(s154,r272,d33,s210,d34);
full_adder fa34(s155,r273,d34,s211,d35);
full_adder fa35(s156,r274,d35,s212,d36);
full_adder fa36(s157,r275,d36,s213,d37);
full_adder fa37(s158,r276,d37,s214,d38);
full_adder fa38(s159,r277,d38,s215,d39);
full_adder fa39(s160,r278,d39,s216,d40);
full_adder fa40(s161,r279,d40,s217,d41);
full_adder fa41(s162,r280,d41,s218,d42);
full_adder fa42(s163,r281,d42,s219,d43);
full_adder fa43(s164,r282,d43,s220,d44);
full_adder fa44(s165,r283,d44,s221,d45);
full_adder fa45(s166,r284,d45,s222,d46);
full_adder fa46(s167,r285,d46,s223,d47);
full_adder fa47(s168,r286,d47,s224,d48);
full_adder fa48(s169,r287,d48,s225,d49);
full_adder fa49(s170,r288,d49,s226,d50);
full_adder fa50(s171,r289,d50,s227,d51);
full_adder fa51(s172,r290,d51,s228,d52);
full_adder fa52(s173,r291,d52,s229,d53);
full_adder fa53(s174,r292,d53,s230,d54);
full_adder fa54(s175,r293,d54,s231,d55);
full_adder fa55(s176,1'b0,d55,s232,d56);
full_adder fa56(s177,1'b0,d56,p61,);

endmodule

module stage4(r294,r295,r296,r297,r298,r299,r300,r301,r302,r303,r304,r305,r306,r307,r308,r309,r310,r311,r312,r313,r314,r315,r316,r317,r318,r319,r320,r321,r322,r323,r324,r325,r326,r327,r328,r329,r330,r331,r332,r333,r334,r335,r336,r337,r338,r339,r340,r341,r342,r343,r344,r345,r346,s178,s179,s180,s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,s226,s227,s228,s229,s230,s231,s232,s233,s234,s235,s236,s237,s238,s239,s240,s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,s256,s257,s258,s259,s260,s261,s262,s263,s264,s265,s266,s267,s268,s269,s270,s271,s272,s273,s274,s275,s276,s277,s278,s279,s280,s281,s282,s283,s284,s285,p6,p60);
input r294,r295,r296,r297,r298,r299,r300,r301,r302,r303,r304,r305,r306,r307,r308,r309,r310,r311,r312,r313,r314,r315,r316,r317,r318,r319,r320,r321,r322,r323,r324,r325,r326,r327,r328,r329,r330,r331,r332,r333,r334,r335,r336,r337,r338,r339,r340,r341,r342,r343,r344,r345,r346,s178,s179,s180,s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,s226,s227,s228,s229,s230,s231,s232;
output s233,s234,s235,s236,s237,s238,s239,s240,s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,s256,s257,s258,s259,s260,s261,s262,s263,s264,s265,s266,s267,s268,s269,s270,s271,s272,s273,s274,s275,s276,s277,s278,s279,s280,s281,s282,s283,s284,s285,p6,p60;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,d49,d50,d51,d52,d53,d54;


full_adder fa0(s178,r294,1'b0,p6,d1);
full_adder fa1(s179,r295,d1,s233,d2);
full_adder fa2(s180,r296,d2,s234,d3);
full_adder fa3(s181,r297,d3,s235,d4);
full_adder fa4(s182,r298,d4,s236,d5);
full_adder fa5(s183,r299,d5,s237,d6);
full_adder fa6(s184,r300,d6,s238,d7);
full_adder fa7(s185,r301,d7,s239,d8);
full_adder fa8(s186,r302,d8,s240,d9);
full_adder fa9(s187,r303,d9,s241,d10);
full_adder fa10(s188,r304,d10,s242,d11);
full_adder fa11(s189,r305,d11,s243,d12);
full_adder fa12(s190,r306,d12,s244,d13);
full_adder fa13(s191,r307,d13,s245,d14);
full_adder fa14(s192,r308,d14,s246,d15);
full_adder fa15(s193,r309,d15,s247,d16);
full_adder fa16(s194,r310,d16,s248,d17);
full_adder fa17(s195,r311,d17,s249,d18);
full_adder fa18(s196,r312,d18,s250,d19);
full_adder fa19(s197,r313,d19,s251,d20);
full_adder fa20(s198,r314,d20,s252,d21);
full_adder fa21(s199,r315,d21,s253,d22);
full_adder fa22(s200,r316,d22,s254,d23);
full_adder fa23(s201,r317,d23,s255,d24);
full_adder fa24(s202,r318,d24,s256,d25);
full_adder fa25(s203,r319,d25,s257,d26);
full_adder fa26(s204,r320,d26,s258,d27);
full_adder fa27(s205,r321,d27,s259,d28);
full_adder fa28(s206,r322,d28,s260,d29);
full_adder fa29(s207,r323,d29,s261,d30);
full_adder fa30(s208,r324,d30,s262,d31);
full_adder fa31(s209,r325,d31,s263,d32);
full_adder fa32(s210,r326,d32,s264,d33);
full_adder fa33(s211,r327,d33,s265,d34);
full_adder fa34(s212,r328,d34,s266,d35);
full_adder fa35(s213,r329,d35,s267,d36);
full_adder fa36(s214,r330,d36,s268,d37);
full_adder fa37(s215,r331,d37,s269,d38);
full_adder fa38(s216,r332,d38,s270,d39);
full_adder fa39(s217,r333,d39,s271,d40);
full_adder fa40(s218,r334,d40,s272,d41);
full_adder fa41(s219,r335,d41,s273,d42);
full_adder fa42(s220,r336,d42,s274,d43);
full_adder fa43(s221,r337,d43,s275,d44);
full_adder fa44(s222,r338,d44,s276,d45);
full_adder fa45(s223,r339,d45,s277,d46);
full_adder fa46(s224,r340,d46,s278,d47);
full_adder fa47(s225,r341,d47,s279,d48);
full_adder fa48(s226,r342,d48,s280,d49);
full_adder fa49(s227,r343,d49,s281,d50);
full_adder fa50(s228,r344,d50,s282,d51);
full_adder fa51(s229,r345,d51,s283,d52);
full_adder fa52(s230,r346,d52,s284,d53);
full_adder fa53(s231,1'b0,d53,s285,d54);
full_adder fa54(s232,1'b0,d54,p60,);

endmodule

module stage5(r347,r348,r349,r350,r351,r352,r353,r354,r355,r356,r357,r358,r359,r360,r361,r362,r363,r364,r365,r366,r367,r368,r369,r370,r371,r372,r373,r374,r375,r376,r377,r378,r379,r380,r381,r382,r383,r384,r385,r386,r387,r388,r389,r390,r391,r392,r393,r394,r395,r396,r397,s233,s234,s235,s236,s237,s238,s239,s240,s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,s256,s257,s258,s259,s260,s261,s262,s263,s264,s265,s266,s267,s268,s269,s270,s271,s272,s273,s274,s275,s276,s277,s278,s279,s280,s281,s282,s283,s284,s285,s286,s287,s288,s289,s290,s291,s292,s293,s294,s295,s296,s297,s298,s299,s300,s301,s302,s303,s304,s305,s306,s307,s308,s309,s310,s311,s312,s313,s314,s315,s316,s317,s318,s319,s320,s321,s322,s323,s324,s325,s326,s327,s328,s329,s330,s331,s332,s333,s334,s335,s336,p7,p59);
input r347,r348,r349,r350,r351,r352,r353,r354,r355,r356,r357,r358,r359,r360,r361,r362,r363,r364,r365,r366,r367,r368,r369,r370,r371,r372,r373,r374,r375,r376,r377,r378,r379,r380,r381,r382,r383,r384,r385,r386,r387,r388,r389,r390,r391,r392,r393,r394,r395,r396,r397,s233,s234,s235,s236,s237,s238,s239,s240,s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,s256,s257,s258,s259,s260,s261,s262,s263,s264,s265,s266,s267,s268,s269,s270,s271,s272,s273,s274,s275,s276,s277,s278,s279,s280,s281,s282,s283,s284,s285;
output s286,s287,s288,s289,s290,s291,s292,s293,s294,s295,s296,s297,s298,s299,s300,s301,s302,s303,s304,s305,s306,s307,s308,s309,s310,s311,s312,s313,s314,s315,s316,s317,s318,s319,s320,s321,s322,s323,s324,s325,s326,s327,s328,s329,s330,s331,s332,s333,s334,s335,s336,p7,p59;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,d49,d50,d51,d52;


full_adder fa0(s233,r347,1'b0,p7,d1);
full_adder fa1(s234,r348,d1,s286,d2);
full_adder fa2(s235,r349,d2,s287,d3);
full_adder fa3(s236,r350,d3,s288,d4);
full_adder fa4(s237,r351,d4,s289,d5);
full_adder fa5(s238,r352,d5,s290,d6);
full_adder fa6(s239,r353,d6,s291,d7);
full_adder fa7(s240,r354,d7,s292,d8);
full_adder fa8(s241,r355,d8,s293,d9);
full_adder fa9(s242,r356,d9,s294,d10);
full_adder fa10(s243,r357,d10,s295,d11);
full_adder fa11(s244,r358,d11,s296,d12);
full_adder fa12(s245,r359,d12,s297,d13);
full_adder fa13(s246,r360,d13,s298,d14);
full_adder fa14(s247,r361,d14,s299,d15);
full_adder fa15(s248,r362,d15,s300,d16);
full_adder fa16(s249,r363,d16,s301,d17);
full_adder fa17(s250,r364,d17,s302,d18);
full_adder fa18(s251,r365,d18,s303,d19);
full_adder fa19(s252,r366,d19,s304,d20);
full_adder fa20(s253,r367,d20,s305,d21);
full_adder fa21(s254,r368,d21,s306,d22);
full_adder fa22(s255,r369,d22,s307,d23);
full_adder fa23(s256,r370,d23,s308,d24);
full_adder fa24(s257,r371,d24,s309,d25);
full_adder fa25(s258,r372,d25,s310,d26);
full_adder fa26(s259,r373,d26,s311,d27);
full_adder fa27(s260,r374,d27,s312,d28);
full_adder fa28(s261,r375,d28,s313,d29);
full_adder fa29(s262,r376,d29,s314,d30);
full_adder fa30(s263,r377,d30,s315,d31);
full_adder fa31(s264,r378,d31,s316,d32);
full_adder fa32(s265,r379,d32,s317,d33);
full_adder fa33(s266,r380,d33,s318,d34);
full_adder fa34(s267,r381,d34,s319,d35);
full_adder fa35(s268,r382,d35,s320,d36);
full_adder fa36(s269,r383,d36,s321,d37);
full_adder fa37(s270,r384,d37,s322,d38);
full_adder fa38(s271,r385,d38,s323,d39);
full_adder fa39(s272,r386,d39,s324,d40);
full_adder fa40(s273,r387,d40,s325,d41);
full_adder fa41(s274,r388,d41,s326,d42);
full_adder fa42(s275,r389,d42,s327,d43);
full_adder fa43(s276,r390,d43,s328,d44);
full_adder fa44(s277,r391,d44,s329,d45);
full_adder fa45(s278,r392,d45,s330,d46);
full_adder fa46(s279,r393,d46,s331,d47);
full_adder fa47(s280,r394,d47,s332,d48);
full_adder fa48(s281,r395,d48,s333,d49);
full_adder fa49(s282,r396,d49,s334,d50);
full_adder fa50(s283,r397,d50,s335,d51);
full_adder fa51(s284,1'b0,d51,s336,d52);
full_adder fa52(s285,1'b0,d52,p59,);

endmodule

module stage6(r398,r399,r400,r401,r402,r403,r404,r405,r406,r407,r408,r409,r410,r411,r412,r413,r414,r415,r416,r417,r418,r419,r420,r421,r422,r423,r424,r425,r426,r427,r428,r429,r430,r431,r432,r433,r434,r435,r436,r437,r438,r439,r440,r441,r442,r443,r444,r445,r446,s286,s287,s288,s289,s290,s291,s292,s293,s294,s295,s296,s297,s298,s299,s300,s301,s302,s303,s304,s305,s306,s307,s308,s309,s310,s311,s312,s313,s314,s315,s316,s317,s318,s319,s320,s321,s322,s323,s324,s325,s326,s327,s328,s329,s330,s331,s332,s333,s334,s335,s336,s337,s338,s339,s340,s341,s342,s343,s344,s345,s346,s347,s348,s349,s350,s351,s352,s353,s354,s355,s356,s357,s358,s359,s360,s361,s362,s363,s364,s365,s366,s367,s368,s369,s370,s371,s372,s373,s374,s375,s376,s377,s378,s379,s380,s381,s382,s383,s384,s385,p8,p58);
input r398,r399,r400,r401,r402,r403,r404,r405,r406,r407,r408,r409,r410,r411,r412,r413,r414,r415,r416,r417,r418,r419,r420,r421,r422,r423,r424,r425,r426,r427,r428,r429,r430,r431,r432,r433,r434,r435,r436,r437,r438,r439,r440,r441,r442,r443,r444,r445,r446,s286,s287,s288,s289,s290,s291,s292,s293,s294,s295,s296,s297,s298,s299,s300,s301,s302,s303,s304,s305,s306,s307,s308,s309,s310,s311,s312,s313,s314,s315,s316,s317,s318,s319,s320,s321,s322,s323,s324,s325,s326,s327,s328,s329,s330,s331,s332,s333,s334,s335,s336;
output s337,s338,s339,s340,s341,s342,s343,s344,s345,s346,s347,s348,s349,s350,s351,s352,s353,s354,s355,s356,s357,s358,s359,s360,s361,s362,s363,s364,s365,s366,s367,s368,s369,s370,s371,s372,s373,s374,s375,s376,s377,s378,s379,s380,s381,s382,s383,s384,s385,p8,p58;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,d49,d50;


full_adder fa0(s286,r398,1'b0,p8,d1);
full_adder fa1(s287,r399,d1,s337,d2);
full_adder fa2(s288,r400,d2,s338,d3);
full_adder fa3(s289,r401,d3,s339,d4);
full_adder fa4(s290,r402,d4,s340,d5);
full_adder fa5(s291,r403,d5,s341,d6);
full_adder fa6(s292,r404,d6,s342,d7);
full_adder fa7(s293,r405,d7,s343,d8);
full_adder fa8(s294,r406,d8,s344,d9);
full_adder fa9(s295,r407,d9,s345,d10);
full_adder fa10(s296,r408,d10,s346,d11);
full_adder fa11(s297,r409,d11,s347,d12);
full_adder fa12(s298,r410,d12,s348,d13);
full_adder fa13(s299,r411,d13,s349,d14);
full_adder fa14(s300,r412,d14,s350,d15);
full_adder fa15(s301,r413,d15,s351,d16);
full_adder fa16(s302,r414,d16,s352,d17);
full_adder fa17(s303,r415,d17,s353,d18);
full_adder fa18(s304,r416,d18,s354,d19);
full_adder fa19(s305,r417,d19,s355,d20);
full_adder fa20(s306,r418,d20,s356,d21);
full_adder fa21(s307,r419,d21,s357,d22);
full_adder fa22(s308,r420,d22,s358,d23);
full_adder fa23(s309,r421,d23,s359,d24);
full_adder fa24(s310,r422,d24,s360,d25);
full_adder fa25(s311,r423,d25,s361,d26);
full_adder fa26(s312,r424,d26,s362,d27);
full_adder fa27(s313,r425,d27,s363,d28);
full_adder fa28(s314,r426,d28,s364,d29);
full_adder fa29(s315,r427,d29,s365,d30);
full_adder fa30(s316,r428,d30,s366,d31);
full_adder fa31(s317,r429,d31,s367,d32);
full_adder fa32(s318,r430,d32,s368,d33);
full_adder fa33(s319,r431,d33,s369,d34);
full_adder fa34(s320,r432,d34,s370,d35);
full_adder fa35(s321,r433,d35,s371,d36);
full_adder fa36(s322,r434,d36,s372,d37);
full_adder fa37(s323,r435,d37,s373,d38);
full_adder fa38(s324,r436,d38,s374,d39);
full_adder fa39(s325,r437,d39,s375,d40);
full_adder fa40(s326,r438,d40,s376,d41);
full_adder fa41(s327,r439,d41,s377,d42);
full_adder fa42(s328,r440,d42,s378,d43);
full_adder fa43(s329,r441,d43,s379,d44);
full_adder fa44(s330,r442,d44,s380,d45);
full_adder fa45(s331,r443,d45,s381,d46);
full_adder fa46(s332,r444,d46,s382,d47);
full_adder fa47(s333,r445,d47,s383,d48);
full_adder fa48(s334,r446,d48,s384,d49);
full_adder fa49(s335,1'b0,d49,s385,d50);
full_adder fa50(s336,1'b0,d50,p58,);

endmodule

module stage7(r447,r448,r449,r450,r451,r452,r453,r454,r455,r456,r457,r458,r459,r460,r461,r462,r463,r464,r465,r466,r467,r468,r469,r470,r471,r472,r473,r474,r475,r476,r477,r478,r479,r480,r481,r482,r483,r484,r485,r486,r487,r488,r489,r490,r491,r492,r493,s337,s338,s339,s340,s341,s342,s343,s344,s345,s346,s347,s348,s349,s350,s351,s352,s353,s354,s355,s356,s357,s358,s359,s360,s361,s362,s363,s364,s365,s366,s367,s368,s369,s370,s371,s372,s373,s374,s375,s376,s377,s378,s379,s380,s381,s382,s383,s384,s385,s386,s387,s388,s389,s390,s391,s392,s393,s394,s395,s396,s397,s398,s399,s400,s401,s402,s403,s404,s405,s406,s407,s408,s409,s410,s411,s412,s413,s414,s415,s416,s417,s418,s419,s420,s421,s422,s423,s424,s425,s426,s427,s428,s429,s430,s431,s432,p9,p57);
input r447,r448,r449,r450,r451,r452,r453,r454,r455,r456,r457,r458,r459,r460,r461,r462,r463,r464,r465,r466,r467,r468,r469,r470,r471,r472,r473,r474,r475,r476,r477,r478,r479,r480,r481,r482,r483,r484,r485,r486,r487,r488,r489,r490,r491,r492,r493,s337,s338,s339,s340,s341,s342,s343,s344,s345,s346,s347,s348,s349,s350,s351,s352,s353,s354,s355,s356,s357,s358,s359,s360,s361,s362,s363,s364,s365,s366,s367,s368,s369,s370,s371,s372,s373,s374,s375,s376,s377,s378,s379,s380,s381,s382,s383,s384,s385;
output s386,s387,s388,s389,s390,s391,s392,s393,s394,s395,s396,s397,s398,s399,s400,s401,s402,s403,s404,s405,s406,s407,s408,s409,s410,s411,s412,s413,s414,s415,s416,s417,s418,s419,s420,s421,s422,s423,s424,s425,s426,s427,s428,s429,s430,s431,s432,p9,p57;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48;


full_adder fa0(s337,r447,1'b0,p9,d1);
full_adder fa1(s338,r448,d1,s386,d2);
full_adder fa2(s339,r449,d2,s387,d3);
full_adder fa3(s340,r450,d3,s388,d4);
full_adder fa4(s341,r451,d4,s389,d5);
full_adder fa5(s342,r452,d5,s390,d6);
full_adder fa6(s343,r453,d6,s391,d7);
full_adder fa7(s344,r454,d7,s392,d8);
full_adder fa8(s345,r455,d8,s393,d9);
full_adder fa9(s346,r456,d9,s394,d10);
full_adder fa10(s347,r457,d10,s395,d11);
full_adder fa11(s348,r458,d11,s396,d12);
full_adder fa12(s349,r459,d12,s397,d13);
full_adder fa13(s350,r460,d13,s398,d14);
full_adder fa14(s351,r461,d14,s399,d15);
full_adder fa15(s352,r462,d15,s400,d16);
full_adder fa16(s353,r463,d16,s401,d17);
full_adder fa17(s354,r464,d17,s402,d18);
full_adder fa18(s355,r465,d18,s403,d19);
full_adder fa19(s356,r466,d19,s404,d20);
full_adder fa20(s357,r467,d20,s405,d21);
full_adder fa21(s358,r468,d21,s406,d22);
full_adder fa22(s359,r469,d22,s407,d23);
full_adder fa23(s360,r470,d23,s408,d24);
full_adder fa24(s361,r471,d24,s409,d25);
full_adder fa25(s362,r472,d25,s410,d26);
full_adder fa26(s363,r473,d26,s411,d27);
full_adder fa27(s364,r474,d27,s412,d28);
full_adder fa28(s365,r475,d28,s413,d29);
full_adder fa29(s366,r476,d29,s414,d30);
full_adder fa30(s367,r477,d30,s415,d31);
full_adder fa31(s368,r478,d31,s416,d32);
full_adder fa32(s369,r479,d32,s417,d33);
full_adder fa33(s370,r480,d33,s418,d34);
full_adder fa34(s371,r481,d34,s419,d35);
full_adder fa35(s372,r482,d35,s420,d36);
full_adder fa36(s373,r483,d36,s421,d37);
full_adder fa37(s374,r484,d37,s422,d38);
full_adder fa38(s375,r485,d38,s423,d39);
full_adder fa39(s376,r486,d39,s424,d40);
full_adder fa40(s377,r487,d40,s425,d41);
full_adder fa41(s378,r488,d41,s426,d42);
full_adder fa42(s379,r489,d42,s427,d43);
full_adder fa43(s380,r490,d43,s428,d44);
full_adder fa44(s381,r491,d44,s429,d45);
full_adder fa45(s382,r492,d45,s430,d46);
full_adder fa46(s383,r493,d46,s431,d47);
full_adder fa47(s384,1'b0,d47,s432,d48);
full_adder fa48(s385,1'b0,d48,p57,);

endmodule

module stage8(r494,r495,r496,r497,r498,r499,r500,r501,r502,r503,r504,r505,r506,r507,r508,r509,r510,r511,r512,r513,r514,r515,r516,r517,r518,r519,r520,r521,r522,r523,r524,r525,r526,r527,r528,r529,r530,r531,r532,r533,r534,r535,r536,r537,r538,s386,s387,s388,s389,s390,s391,s392,s393,s394,s395,s396,s397,s398,s399,s400,s401,s402,s403,s404,s405,s406,s407,s408,s409,s410,s411,s412,s413,s414,s415,s416,s417,s418,s419,s420,s421,s422,s423,s424,s425,s426,s427,s428,s429,s430,s431,s432,s433,s434,s435,s436,s437,s438,s439,s440,s441,s442,s443,s444,s445,s446,s447,s448,s449,s450,s451,s452,s453,s454,s455,s456,s457,s458,s459,s460,s461,s462,s463,s464,s465,s466,s467,s468,s469,s470,s471,s472,s473,s474,s475,s476,s477,p10,p56);
input r494,r495,r496,r497,r498,r499,r500,r501,r502,r503,r504,r505,r506,r507,r508,r509,r510,r511,r512,r513,r514,r515,r516,r517,r518,r519,r520,r521,r522,r523,r524,r525,r526,r527,r528,r529,r530,r531,r532,r533,r534,r535,r536,r537,r538,s386,s387,s388,s389,s390,s391,s392,s393,s394,s395,s396,s397,s398,s399,s400,s401,s402,s403,s404,s405,s406,s407,s408,s409,s410,s411,s412,s413,s414,s415,s416,s417,s418,s419,s420,s421,s422,s423,s424,s425,s426,s427,s428,s429,s430,s431,s432;
output s433,s434,s435,s436,s437,s438,s439,s440,s441,s442,s443,s444,s445,s446,s447,s448,s449,s450,s451,s452,s453,s454,s455,s456,s457,s458,s459,s460,s461,s462,s463,s464,s465,s466,s467,s468,s469,s470,s471,s472,s473,s474,s475,s476,s477,p10,p56;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46;


full_adder fa0(s386,r494,1'b0,p10,d1);
full_adder fa1(s387,r495,d1,s433,d2);
full_adder fa2(s388,r496,d2,s434,d3);
full_adder fa3(s389,r497,d3,s435,d4);
full_adder fa4(s390,r498,d4,s436,d5);
full_adder fa5(s391,r499,d5,s437,d6);
full_adder fa6(s392,r500,d6,s438,d7);
full_adder fa7(s393,r501,d7,s439,d8);
full_adder fa8(s394,r502,d8,s440,d9);
full_adder fa9(s395,r503,d9,s441,d10);
full_adder fa10(s396,r504,d10,s442,d11);
full_adder fa11(s397,r505,d11,s443,d12);
full_adder fa12(s398,r506,d12,s444,d13);
full_adder fa13(s399,r507,d13,s445,d14);
full_adder fa14(s400,r508,d14,s446,d15);
full_adder fa15(s401,r509,d15,s447,d16);
full_adder fa16(s402,r510,d16,s448,d17);
full_adder fa17(s403,r511,d17,s449,d18);
full_adder fa18(s404,r512,d18,s450,d19);
full_adder fa19(s405,r513,d19,s451,d20);
full_adder fa20(s406,r514,d20,s452,d21);
full_adder fa21(s407,r515,d21,s453,d22);
full_adder fa22(s408,r516,d22,s454,d23);
full_adder fa23(s409,r517,d23,s455,d24);
full_adder fa24(s410,r518,d24,s456,d25);
full_adder fa25(s411,r519,d25,s457,d26);
full_adder fa26(s412,r520,d26,s458,d27);
full_adder fa27(s413,r521,d27,s459,d28);
full_adder fa28(s414,r522,d28,s460,d29);
full_adder fa29(s415,r523,d29,s461,d30);
full_adder fa30(s416,r524,d30,s462,d31);
full_adder fa31(s417,r525,d31,s463,d32);
full_adder fa32(s418,r526,d32,s464,d33);
full_adder fa33(s419,r527,d33,s465,d34);
full_adder fa34(s420,r528,d34,s466,d35);
full_adder fa35(s421,r529,d35,s467,d36);
full_adder fa36(s422,r530,d36,s468,d37);
full_adder fa37(s423,r531,d37,s469,d38);
full_adder fa38(s424,r532,d38,s470,d39);
full_adder fa39(s425,r533,d39,s471,d40);
full_adder fa40(s426,r534,d40,s472,d41);
full_adder fa41(s427,r535,d41,s473,d42);
full_adder fa42(s428,r536,d42,s474,d43);
full_adder fa43(s429,r537,d43,s475,d44);
full_adder fa44(s430,r538,d44,s476,d45);
full_adder fa45(s431,1'b0,d45,s477,d46);
full_adder fa46(s432,1'b0,d46,p56,);

endmodule

module stage9(r539,r540,r541,r542,r543,r544,r545,r546,r547,r548,r549,r550,r551,r552,r553,r554,r555,r556,r557,r558,r559,r560,r561,r562,r563,r564,r565,r566,r567,r568,r569,r570,r571,r572,r573,r574,r575,r576,r577,r578,r579,r580,r581,s433,s434,s435,s436,s437,s438,s439,s440,s441,s442,s443,s444,s445,s446,s447,s448,s449,s450,s451,s452,s453,s454,s455,s456,s457,s458,s459,s460,s461,s462,s463,s464,s465,s466,s467,s468,s469,s470,s471,s472,s473,s474,s475,s476,s477,s478,s479,s480,s481,s482,s483,s484,s485,s486,s487,s488,s489,s490,s491,s492,s493,s494,s495,s496,s497,s498,s499,s500,s501,s502,s503,s504,s505,s506,s507,s508,s509,s510,s511,s512,s513,s514,s515,s516,s517,s518,s519,s520,p11,p55);
input r539,r540,r541,r542,r543,r544,r545,r546,r547,r548,r549,r550,r551,r552,r553,r554,r555,r556,r557,r558,r559,r560,r561,r562,r563,r564,r565,r566,r567,r568,r569,r570,r571,r572,r573,r574,r575,r576,r577,r578,r579,r580,r581,s433,s434,s435,s436,s437,s438,s439,s440,s441,s442,s443,s444,s445,s446,s447,s448,s449,s450,s451,s452,s453,s454,s455,s456,s457,s458,s459,s460,s461,s462,s463,s464,s465,s466,s467,s468,s469,s470,s471,s472,s473,s474,s475,s476,s477;
output s478,s479,s480,s481,s482,s483,s484,s485,s486,s487,s488,s489,s490,s491,s492,s493,s494,s495,s496,s497,s498,s499,s500,s501,s502,s503,s504,s505,s506,s507,s508,s509,s510,s511,s512,s513,s514,s515,s516,s517,s518,s519,s520,p11,p55;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44;


full_adder fa0(s433,r539,1'b0,p11,d1);
full_adder fa1(s434,r540,d1,s478,d2);
full_adder fa2(s435,r541,d2,s479,d3);
full_adder fa3(s436,r542,d3,s480,d4);
full_adder fa4(s437,r543,d4,s481,d5);
full_adder fa5(s438,r544,d5,s482,d6);
full_adder fa6(s439,r545,d6,s483,d7);
full_adder fa7(s440,r546,d7,s484,d8);
full_adder fa8(s441,r547,d8,s485,d9);
full_adder fa9(s442,r548,d9,s486,d10);
full_adder fa10(s443,r549,d10,s487,d11);
full_adder fa11(s444,r550,d11,s488,d12);
full_adder fa12(s445,r551,d12,s489,d13);
full_adder fa13(s446,r552,d13,s490,d14);
full_adder fa14(s447,r553,d14,s491,d15);
full_adder fa15(s448,r554,d15,s492,d16);
full_adder fa16(s449,r555,d16,s493,d17);
full_adder fa17(s450,r556,d17,s494,d18);
full_adder fa18(s451,r557,d18,s495,d19);
full_adder fa19(s452,r558,d19,s496,d20);
full_adder fa20(s453,r559,d20,s497,d21);
full_adder fa21(s454,r560,d21,s498,d22);
full_adder fa22(s455,r561,d22,s499,d23);
full_adder fa23(s456,r562,d23,s500,d24);
full_adder fa24(s457,r563,d24,s501,d25);
full_adder fa25(s458,r564,d25,s502,d26);
full_adder fa26(s459,r565,d26,s503,d27);
full_adder fa27(s460,r566,d27,s504,d28);
full_adder fa28(s461,r567,d28,s505,d29);
full_adder fa29(s462,r568,d29,s506,d30);
full_adder fa30(s463,r569,d30,s507,d31);
full_adder fa31(s464,r570,d31,s508,d32);
full_adder fa32(s465,r571,d32,s509,d33);
full_adder fa33(s466,r572,d33,s510,d34);
full_adder fa34(s467,r573,d34,s511,d35);
full_adder fa35(s468,r574,d35,s512,d36);
full_adder fa36(s469,r575,d36,s513,d37);
full_adder fa37(s470,r576,d37,s514,d38);
full_adder fa38(s471,r577,d38,s515,d39);
full_adder fa39(s472,r578,d39,s516,d40);
full_adder fa40(s473,r579,d40,s517,d41);
full_adder fa41(s474,r580,d41,s518,d42);
full_adder fa42(s475,r581,d42,s519,d43);
full_adder fa43(s476,1'b0,d43,s520,d44);
full_adder fa44(s477,1'b0,d44,p55,);

endmodule

module stage10(r582,r583,r584,r585,r586,r587,r588,r589,r590,r591,r592,r593,r594,r595,r596,r597,r598,r599,r600,r601,r602,r603,r604,r605,r606,r607,r608,r609,r610,r611,r612,r613,r614,r615,r616,r617,r618,r619,r620,r621,r622,s478,s479,s480,s481,s482,s483,s484,s485,s486,s487,s488,s489,s490,s491,s492,s493,s494,s495,s496,s497,s498,s499,s500,s501,s502,s503,s504,s505,s506,s507,s508,s509,s510,s511,s512,s513,s514,s515,s516,s517,s518,s519,s520,s521,s522,s523,s524,s525,s526,s527,s528,s529,s530,s531,s532,s533,s534,s535,s536,s537,s538,s539,s540,s541,s542,s543,s544,s545,s546,s547,s548,s549,s550,s551,s552,s553,s554,s555,s556,s557,s558,s559,s560,s561,p12,p54);
input r582,r583,r584,r585,r586,r587,r588,r589,r590,r591,r592,r593,r594,r595,r596,r597,r598,r599,r600,r601,r602,r603,r604,r605,r606,r607,r608,r609,r610,r611,r612,r613,r614,r615,r616,r617,r618,r619,r620,r621,r622,s478,s479,s480,s481,s482,s483,s484,s485,s486,s487,s488,s489,s490,s491,s492,s493,s494,s495,s496,s497,s498,s499,s500,s501,s502,s503,s504,s505,s506,s507,s508,s509,s510,s511,s512,s513,s514,s515,s516,s517,s518,s519,s520;
output s521,s522,s523,s524,s525,s526,s527,s528,s529,s530,s531,s532,s533,s534,s535,s536,s537,s538,s539,s540,s541,s542,s543,s544,s545,s546,s547,s548,s549,s550,s551,s552,s553,s554,s555,s556,s557,s558,s559,s560,s561,p12,p54;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42;


full_adder fa0(s478,r582,1'b0,p12,d1);
full_adder fa1(s479,r583,d1,s521,d2);
full_adder fa2(s480,r584,d2,s522,d3);
full_adder fa3(s481,r585,d3,s523,d4);
full_adder fa4(s482,r586,d4,s524,d5);
full_adder fa5(s483,r587,d5,s525,d6);
full_adder fa6(s484,r588,d6,s526,d7);
full_adder fa7(s485,r589,d7,s527,d8);
full_adder fa8(s486,r590,d8,s528,d9);
full_adder fa9(s487,r591,d9,s529,d10);
full_adder fa10(s488,r592,d10,s530,d11);
full_adder fa11(s489,r593,d11,s531,d12);
full_adder fa12(s490,r594,d12,s532,d13);
full_adder fa13(s491,r595,d13,s533,d14);
full_adder fa14(s492,r596,d14,s534,d15);
full_adder fa15(s493,r597,d15,s535,d16);
full_adder fa16(s494,r598,d16,s536,d17);
full_adder fa17(s495,r599,d17,s537,d18);
full_adder fa18(s496,r600,d18,s538,d19);
full_adder fa19(s497,r601,d19,s539,d20);
full_adder fa20(s498,r602,d20,s540,d21);
full_adder fa21(s499,r603,d21,s541,d22);
full_adder fa22(s500,r604,d22,s542,d23);
full_adder fa23(s501,r605,d23,s543,d24);
full_adder fa24(s502,r606,d24,s544,d25);
full_adder fa25(s503,r607,d25,s545,d26);
full_adder fa26(s504,r608,d26,s546,d27);
full_adder fa27(s505,r609,d27,s547,d28);
full_adder fa28(s506,r610,d28,s548,d29);
full_adder fa29(s507,r611,d29,s549,d30);
full_adder fa30(s508,r612,d30,s550,d31);
full_adder fa31(s509,r613,d31,s551,d32);
full_adder fa32(s510,r614,d32,s552,d33);
full_adder fa33(s511,r615,d33,s553,d34);
full_adder fa34(s512,r616,d34,s554,d35);
full_adder fa35(s513,r617,d35,s555,d36);
full_adder fa36(s514,r618,d36,s556,d37);
full_adder fa37(s515,r619,d37,s557,d38);
full_adder fa38(s516,r620,d38,s558,d39);
full_adder fa39(s517,r621,d39,s559,d40);
full_adder fa40(s518,r622,d40,s560,d41);
full_adder fa41(s519,1'b0,d41,s561,d42);
full_adder fa42(s520,1'b0,d42,p54,);

endmodule

module stage11(r623,r624,r625,r626,r627,r628,r629,r630,r631,r632,r633,r634,r635,r636,r637,r638,r639,r640,r641,r642,r643,r644,r645,r646,r647,r648,r649,r650,r651,r652,r653,r654,r655,r656,r657,r658,r659,r660,r661,s521,s522,s523,s524,s525,s526,s527,s528,s529,s530,s531,s532,s533,s534,s535,s536,s537,s538,s539,s540,s541,s542,s543,s544,s545,s546,s547,s548,s549,s550,s551,s552,s553,s554,s555,s556,s557,s558,s559,s560,s561,s562,s563,s564,s565,s566,s567,s568,s569,s570,s571,s572,s573,s574,s575,s576,s577,s578,s579,s580,s581,s582,s583,s584,s585,s586,s587,s588,s589,s590,s591,s592,s593,s594,s595,s596,s597,s598,s599,s600,p13,p53);
input r623,r624,r625,r626,r627,r628,r629,r630,r631,r632,r633,r634,r635,r636,r637,r638,r639,r640,r641,r642,r643,r644,r645,r646,r647,r648,r649,r650,r651,r652,r653,r654,r655,r656,r657,r658,r659,r660,r661,s521,s522,s523,s524,s525,s526,s527,s528,s529,s530,s531,s532,s533,s534,s535,s536,s537,s538,s539,s540,s541,s542,s543,s544,s545,s546,s547,s548,s549,s550,s551,s552,s553,s554,s555,s556,s557,s558,s559,s560,s561;
output s562,s563,s564,s565,s566,s567,s568,s569,s570,s571,s572,s573,s574,s575,s576,s577,s578,s579,s580,s581,s582,s583,s584,s585,s586,s587,s588,s589,s590,s591,s592,s593,s594,s595,s596,s597,s598,s599,s600,p13,p53;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40;


full_adder fa0(s521,r623,1'b0,p13,d1);
full_adder fa1(s522,r624,d1,s562,d2);
full_adder fa2(s523,r625,d2,s563,d3);
full_adder fa3(s524,r626,d3,s564,d4);
full_adder fa4(s525,r627,d4,s565,d5);
full_adder fa5(s526,r628,d5,s566,d6);
full_adder fa6(s527,r629,d6,s567,d7);
full_adder fa7(s528,r630,d7,s568,d8);
full_adder fa8(s529,r631,d8,s569,d9);
full_adder fa9(s530,r632,d9,s570,d10);
full_adder fa10(s531,r633,d10,s571,d11);
full_adder fa11(s532,r634,d11,s572,d12);
full_adder fa12(s533,r635,d12,s573,d13);
full_adder fa13(s534,r636,d13,s574,d14);
full_adder fa14(s535,r637,d14,s575,d15);
full_adder fa15(s536,r638,d15,s576,d16);
full_adder fa16(s537,r639,d16,s577,d17);
full_adder fa17(s538,r640,d17,s578,d18);
full_adder fa18(s539,r641,d18,s579,d19);
full_adder fa19(s540,r642,d19,s580,d20);
full_adder fa20(s541,r643,d20,s581,d21);
full_adder fa21(s542,r644,d21,s582,d22);
full_adder fa22(s543,r645,d22,s583,d23);
full_adder fa23(s544,r646,d23,s584,d24);
full_adder fa24(s545,r647,d24,s585,d25);
full_adder fa25(s546,r648,d25,s586,d26);
full_adder fa26(s547,r649,d26,s587,d27);
full_adder fa27(s548,r650,d27,s588,d28);
full_adder fa28(s549,r651,d28,s589,d29);
full_adder fa29(s550,r652,d29,s590,d30);
full_adder fa30(s551,r653,d30,s591,d31);
full_adder fa31(s552,r654,d31,s592,d32);
full_adder fa32(s553,r655,d32,s593,d33);
full_adder fa33(s554,r656,d33,s594,d34);
full_adder fa34(s555,r657,d34,s595,d35);
full_adder fa35(s556,r658,d35,s596,d36);
full_adder fa36(s557,r659,d36,s597,d37);
full_adder fa37(s558,r660,d37,s598,d38);
full_adder fa38(s559,r661,d38,s599,d39);
full_adder fa39(s560,1'b0,d39,s600,d40);
full_adder fa40(s561,1'b0,d40,p53,);

endmodule

module stage12(r662,r663,r664,r665,r666,r667,r668,r669,r670,r671,r672,r673,r674,r675,r676,r677,r678,r679,r680,r681,r682,r683,r684,r685,r686,r687,r688,r689,r690,r691,r692,r693,r694,r695,r696,r697,r698,s562,s563,s564,s565,s566,s567,s568,s569,s570,s571,s572,s573,s574,s575,s576,s577,s578,s579,s580,s581,s582,s583,s584,s585,s586,s587,s588,s589,s590,s591,s592,s593,s594,s595,s596,s597,s598,s599,s600,s601,s602,s603,s604,s605,s606,s607,s608,s609,s610,s611,s612,s613,s614,s615,s616,s617,s618,s619,s620,s621,s622,s623,s624,s625,s626,s627,s628,s629,s630,s631,s632,s633,s634,s635,s636,s637,p14,p52);
input r662,r663,r664,r665,r666,r667,r668,r669,r670,r671,r672,r673,r674,r675,r676,r677,r678,r679,r680,r681,r682,r683,r684,r685,r686,r687,r688,r689,r690,r691,r692,r693,r694,r695,r696,r697,r698,s562,s563,s564,s565,s566,s567,s568,s569,s570,s571,s572,s573,s574,s575,s576,s577,s578,s579,s580,s581,s582,s583,s584,s585,s586,s587,s588,s589,s590,s591,s592,s593,s594,s595,s596,s597,s598,s599,s600;
output s601,s602,s603,s604,s605,s606,s607,s608,s609,s610,s611,s612,s613,s614,s615,s616,s617,s618,s619,s620,s621,s622,s623,s624,s625,s626,s627,s628,s629,s630,s631,s632,s633,s634,s635,s636,s637,p14,p52;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38;


full_adder fa0(s562,r662,1'b0,p14,d1);
full_adder fa1(s563,r663,d1,s601,d2);
full_adder fa2(s564,r664,d2,s602,d3);
full_adder fa3(s565,r665,d3,s603,d4);
full_adder fa4(s566,r666,d4,s604,d5);
full_adder fa5(s567,r667,d5,s605,d6);
full_adder fa6(s568,r668,d6,s606,d7);
full_adder fa7(s569,r669,d7,s607,d8);
full_adder fa8(s570,r670,d8,s608,d9);
full_adder fa9(s571,r671,d9,s609,d10);
full_adder fa10(s572,r672,d10,s610,d11);
full_adder fa11(s573,r673,d11,s611,d12);
full_adder fa12(s574,r674,d12,s612,d13);
full_adder fa13(s575,r675,d13,s613,d14);
full_adder fa14(s576,r676,d14,s614,d15);
full_adder fa15(s577,r677,d15,s615,d16);
full_adder fa16(s578,r678,d16,s616,d17);
full_adder fa17(s579,r679,d17,s617,d18);
full_adder fa18(s580,r680,d18,s618,d19);
full_adder fa19(s581,r681,d19,s619,d20);
full_adder fa20(s582,r682,d20,s620,d21);
full_adder fa21(s583,r683,d21,s621,d22);
full_adder fa22(s584,r684,d22,s622,d23);
full_adder fa23(s585,r685,d23,s623,d24);
full_adder fa24(s586,r686,d24,s624,d25);
full_adder fa25(s587,r687,d25,s625,d26);
full_adder fa26(s588,r688,d26,s626,d27);
full_adder fa27(s589,r689,d27,s627,d28);
full_adder fa28(s590,r690,d28,s628,d29);
full_adder fa29(s591,r691,d29,s629,d30);
full_adder fa30(s592,r692,d30,s630,d31);
full_adder fa31(s593,r693,d31,s631,d32);
full_adder fa32(s594,r694,d32,s632,d33);
full_adder fa33(s595,r695,d33,s633,d34);
full_adder fa34(s596,r696,d34,s634,d35);
full_adder fa35(s597,r697,d35,s635,d36);
full_adder fa36(s598,r698,d36,s636,d37);
full_adder fa37(s599,1'b0,d37,s637,d38);
full_adder fa38(s600,1'b0,d38,p52,);

endmodule

module stage13(r699,r700,r701,r702,r703,r704,r705,r706,r707,r708,r709,r710,r711,r712,r713,r714,r715,r716,r717,r718,r719,r720,r721,r722,r723,r724,r725,r726,r727,r728,r729,r730,r731,r732,r733,s601,s602,s603,s604,s605,s606,s607,s608,s609,s610,s611,s612,s613,s614,s615,s616,s617,s618,s619,s620,s621,s622,s623,s624,s625,s626,s627,s628,s629,s630,s631,s632,s633,s634,s635,s636,s637,s638,s639,s640,s641,s642,s643,s644,s645,s646,s647,s648,s649,s650,s651,s652,s653,s654,s655,s656,s657,s658,s659,s660,s661,s662,s663,s664,s665,s666,s667,s668,s669,s670,s671,s672,p15,p51);
input r699,r700,r701,r702,r703,r704,r705,r706,r707,r708,r709,r710,r711,r712,r713,r714,r715,r716,r717,r718,r719,r720,r721,r722,r723,r724,r725,r726,r727,r728,r729,r730,r731,r732,r733,s601,s602,s603,s604,s605,s606,s607,s608,s609,s610,s611,s612,s613,s614,s615,s616,s617,s618,s619,s620,s621,s622,s623,s624,s625,s626,s627,s628,s629,s630,s631,s632,s633,s634,s635,s636,s637;
output s638,s639,s640,s641,s642,s643,s644,s645,s646,s647,s648,s649,s650,s651,s652,s653,s654,s655,s656,s657,s658,s659,s660,s661,s662,s663,s664,s665,s666,s667,s668,s669,s670,s671,s672,p15,p51;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36;


full_adder fa0(s601,r699,1'b0,p15,d1);
full_adder fa1(s602,r700,d1,s638,d2);
full_adder fa2(s603,r701,d2,s639,d3);
full_adder fa3(s604,r702,d3,s640,d4);
full_adder fa4(s605,r703,d4,s641,d5);
full_adder fa5(s606,r704,d5,s642,d6);
full_adder fa6(s607,r705,d6,s643,d7);
full_adder fa7(s608,r706,d7,s644,d8);
full_adder fa8(s609,r707,d8,s645,d9);
full_adder fa9(s610,r708,d9,s646,d10);
full_adder fa10(s611,r709,d10,s647,d11);
full_adder fa11(s612,r710,d11,s648,d12);
full_adder fa12(s613,r711,d12,s649,d13);
full_adder fa13(s614,r712,d13,s650,d14);
full_adder fa14(s615,r713,d14,s651,d15);
full_adder fa15(s616,r714,d15,s652,d16);
full_adder fa16(s617,r715,d16,s653,d17);
full_adder fa17(s618,r716,d17,s654,d18);
full_adder fa18(s619,r717,d18,s655,d19);
full_adder fa19(s620,r718,d19,s656,d20);
full_adder fa20(s621,r719,d20,s657,d21);
full_adder fa21(s622,r720,d21,s658,d22);
full_adder fa22(s623,r721,d22,s659,d23);
full_adder fa23(s624,r722,d23,s660,d24);
full_adder fa24(s625,r723,d24,s661,d25);
full_adder fa25(s626,r724,d25,s662,d26);
full_adder fa26(s627,r725,d26,s663,d27);
full_adder fa27(s628,r726,d27,s664,d28);
full_adder fa28(s629,r727,d28,s665,d29);
full_adder fa29(s630,r728,d29,s666,d30);
full_adder fa30(s631,r729,d30,s667,d31);
full_adder fa31(s632,r730,d31,s668,d32);
full_adder fa32(s633,r731,d32,s669,d33);
full_adder fa33(s634,r732,d33,s670,d34);
full_adder fa34(s635,r733,d34,s671,d35);
full_adder fa35(s636,1'b0,d35,s672,d36);
full_adder fa36(s637,1'b0,d36,p51,);

endmodule

module stage14(r734,r735,r736,r737,r738,r739,r740,r741,r742,r743,r744,r745,r746,r747,r748,r749,r750,r751,r752,r753,r754,r755,r756,r757,r758,r759,r760,r761,r762,r763,r764,r765,r766,s638,s639,s640,s641,s642,s643,s644,s645,s646,s647,s648,s649,s650,s651,s652,s653,s654,s655,s656,s657,s658,s659,s660,s661,s662,s663,s664,s665,s666,s667,s668,s669,s670,s671,s672,s673,s674,s675,s676,s677,s678,s679,s680,s681,s682,s683,s684,s685,s686,s687,s688,s689,s690,s691,s692,s693,s694,s695,s696,s697,s698,s699,s700,s701,s702,s703,s704,s705,p16,p50);
input r734,r735,r736,r737,r738,r739,r740,r741,r742,r743,r744,r745,r746,r747,r748,r749,r750,r751,r752,r753,r754,r755,r756,r757,r758,r759,r760,r761,r762,r763,r764,r765,r766,s638,s639,s640,s641,s642,s643,s644,s645,s646,s647,s648,s649,s650,s651,s652,s653,s654,s655,s656,s657,s658,s659,s660,s661,s662,s663,s664,s665,s666,s667,s668,s669,s670,s671,s672;
output s673,s674,s675,s676,s677,s678,s679,s680,s681,s682,s683,s684,s685,s686,s687,s688,s689,s690,s691,s692,s693,s694,s695,s696,s697,s698,s699,s700,s701,s702,s703,s704,s705,p16,p50;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34;


full_adder fa0(s638,r734,1'b0,p16,d1);
full_adder fa1(s639,r735,d1,s673,d2);
full_adder fa2(s640,r736,d2,s674,d3);
full_adder fa3(s641,r737,d3,s675,d4);
full_adder fa4(s642,r738,d4,s676,d5);
full_adder fa5(s643,r739,d5,s677,d6);
full_adder fa6(s644,r740,d6,s678,d7);
full_adder fa7(s645,r741,d7,s679,d8);
full_adder fa8(s646,r742,d8,s680,d9);
full_adder fa9(s647,r743,d9,s681,d10);
full_adder fa10(s648,r744,d10,s682,d11);
full_adder fa11(s649,r745,d11,s683,d12);
full_adder fa12(s650,r746,d12,s684,d13);
full_adder fa13(s651,r747,d13,s685,d14);
full_adder fa14(s652,r748,d14,s686,d15);
full_adder fa15(s653,r749,d15,s687,d16);
full_adder fa16(s654,r750,d16,s688,d17);
full_adder fa17(s655,r751,d17,s689,d18);
full_adder fa18(s656,r752,d18,s690,d19);
full_adder fa19(s657,r753,d19,s691,d20);
full_adder fa20(s658,r754,d20,s692,d21);
full_adder fa21(s659,r755,d21,s693,d22);
full_adder fa22(s660,r756,d22,s694,d23);
full_adder fa23(s661,r757,d23,s695,d24);
full_adder fa24(s662,r758,d24,s696,d25);
full_adder fa25(s663,r759,d25,s697,d26);
full_adder fa26(s664,r760,d26,s698,d27);
full_adder fa27(s665,r761,d27,s699,d28);
full_adder fa28(s666,r762,d28,s700,d29);
full_adder fa29(s667,r763,d29,s701,d30);
full_adder fa30(s668,r764,d30,s702,d31);
full_adder fa31(s669,r765,d31,s703,d32);
full_adder fa32(s670,r766,d32,s704,d33);
full_adder fa33(s671,1'b0,d33,s705,d34);
full_adder fa34(s672,1'b0,d34,p50,);

endmodule

module stage15(r767,r768,r769,r770,r771,r772,r773,r774,r775,r776,r777,r778,r779,r780,r781,r782,r783,r784,r785,r786,r787,r788,r789,r790,r791,r792,r793,r794,r795,r796,r797,s673,s674,s675,s676,s677,s678,s679,s680,s681,s682,s683,s684,s685,s686,s687,s688,s689,s690,s691,s692,s693,s694,s695,s696,s697,s698,s699,s700,s701,s702,s703,s704,s705,s706,s707,s708,s709,s710,s711,s712,s713,s714,s715,s716,s717,s718,s719,s720,s721,s722,s723,s724,s725,s726,s727,s728,s729,s730,s731,s732,s733,s734,s735,s736,p17,p49);
input r767,r768,r769,r770,r771,r772,r773,r774,r775,r776,r777,r778,r779,r780,r781,r782,r783,r784,r785,r786,r787,r788,r789,r790,r791,r792,r793,r794,r795,r796,r797,s673,s674,s675,s676,s677,s678,s679,s680,s681,s682,s683,s684,s685,s686,s687,s688,s689,s690,s691,s692,s693,s694,s695,s696,s697,s698,s699,s700,s701,s702,s703,s704,s705;
output s706,s707,s708,s709,s710,s711,s712,s713,s714,s715,s716,s717,s718,s719,s720,s721,s722,s723,s724,s725,s726,s727,s728,s729,s730,s731,s732,s733,s734,s735,s736,p17,p49;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32;


full_adder fa0(s673,r767,1'b0,p17,d1);
full_adder fa1(s674,r768,d1,s706,d2);
full_adder fa2(s675,r769,d2,s707,d3);
full_adder fa3(s676,r770,d3,s708,d4);
full_adder fa4(s677,r771,d4,s709,d5);
full_adder fa5(s678,r772,d5,s710,d6);
full_adder fa6(s679,r773,d6,s711,d7);
full_adder fa7(s680,r774,d7,s712,d8);
full_adder fa8(s681,r775,d8,s713,d9);
full_adder fa9(s682,r776,d9,s714,d10);
full_adder fa10(s683,r777,d10,s715,d11);
full_adder fa11(s684,r778,d11,s716,d12);
full_adder fa12(s685,r779,d12,s717,d13);
full_adder fa13(s686,r780,d13,s718,d14);
full_adder fa14(s687,r781,d14,s719,d15);
full_adder fa15(s688,r782,d15,s720,d16);
full_adder fa16(s689,r783,d16,s721,d17);
full_adder fa17(s690,r784,d17,s722,d18);
full_adder fa18(s691,r785,d18,s723,d19);
full_adder fa19(s692,r786,d19,s724,d20);
full_adder fa20(s693,r787,d20,s725,d21);
full_adder fa21(s694,r788,d21,s726,d22);
full_adder fa22(s695,r789,d22,s727,d23);
full_adder fa23(s696,r790,d23,s728,d24);
full_adder fa24(s697,r791,d24,s729,d25);
full_adder fa25(s698,r792,d25,s730,d26);
full_adder fa26(s699,r793,d26,s731,d27);
full_adder fa27(s700,r794,d27,s732,d28);
full_adder fa28(s701,r795,d28,s733,d29);
full_adder fa29(s702,r796,d29,s734,d30);
full_adder fa30(s703,r797,d30,s735,d31);
full_adder fa31(s704,1'b0,d31,s736,d32);
full_adder fa32(s705,1'b0,d32,p49,);

endmodule

module stage16(r798,r799,r800,r801,r802,r803,r804,r805,r806,r807,r808,r809,r810,r811,r812,r813,r814,r815,r816,r817,r818,r819,r820,r821,r822,r823,r824,r825,r826,s706,s707,s708,s709,s710,s711,s712,s713,s714,s715,s716,s717,s718,s719,s720,s721,s722,s723,s724,s725,s726,s727,s728,s729,s730,s731,s732,s733,s734,s735,s736,s737,s738,s739,s740,s741,s742,s743,s744,s745,s746,s747,s748,s749,s750,s751,s752,s753,s754,s755,s756,s757,s758,s759,s760,s761,s762,s763,s764,s765,p18,p48);
input r798,r799,r800,r801,r802,r803,r804,r805,r806,r807,r808,r809,r810,r811,r812,r813,r814,r815,r816,r817,r818,r819,r820,r821,r822,r823,r824,r825,r826,s706,s707,s708,s709,s710,s711,s712,s713,s714,s715,s716,s717,s718,s719,s720,s721,s722,s723,s724,s725,s726,s727,s728,s729,s730,s731,s732,s733,s734,s735,s736;
output s737,s738,s739,s740,s741,s742,s743,s744,s745,s746,s747,s748,s749,s750,s751,s752,s753,s754,s755,s756,s757,s758,s759,s760,s761,s762,s763,s764,s765,p18,p48;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30;


full_adder fa0(s706,r798,1'b0,p18,d1);
full_adder fa1(s707,r799,d1,s737,d2);
full_adder fa2(s708,r800,d2,s738,d3);
full_adder fa3(s709,r801,d3,s739,d4);
full_adder fa4(s710,r802,d4,s740,d5);
full_adder fa5(s711,r803,d5,s741,d6);
full_adder fa6(s712,r804,d6,s742,d7);
full_adder fa7(s713,r805,d7,s743,d8);
full_adder fa8(s714,r806,d8,s744,d9);
full_adder fa9(s715,r807,d9,s745,d10);
full_adder fa10(s716,r808,d10,s746,d11);
full_adder fa11(s717,r809,d11,s747,d12);
full_adder fa12(s718,r810,d12,s748,d13);
full_adder fa13(s719,r811,d13,s749,d14);
full_adder fa14(s720,r812,d14,s750,d15);
full_adder fa15(s721,r813,d15,s751,d16);
full_adder fa16(s722,r814,d16,s752,d17);
full_adder fa17(s723,r815,d17,s753,d18);
full_adder fa18(s724,r816,d18,s754,d19);
full_adder fa19(s725,r817,d19,s755,d20);
full_adder fa20(s726,r818,d20,s756,d21);
full_adder fa21(s727,r819,d21,s757,d22);
full_adder fa22(s728,r820,d22,s758,d23);
full_adder fa23(s729,r821,d23,s759,d24);
full_adder fa24(s730,r822,d24,s760,d25);
full_adder fa25(s731,r823,d25,s761,d26);
full_adder fa26(s732,r824,d26,s762,d27);
full_adder fa27(s733,r825,d27,s763,d28);
full_adder fa28(s734,r826,d28,s764,d29);
full_adder fa29(s735,1'b0,d29,s765,d30);
full_adder fa30(s736,1'b0,d30,p48,);

endmodule

module stage17(r827,r828,r829,r830,r831,r832,r833,r834,r835,r836,r837,r838,r839,r840,r841,r842,r843,r844,r845,r846,r847,r848,r849,r850,r851,r852,r853,s737,s738,s739,s740,s741,s742,s743,s744,s745,s746,s747,s748,s749,s750,s751,s752,s753,s754,s755,s756,s757,s758,s759,s760,s761,s762,s763,s764,s765,s766,s767,s768,s769,s770,s771,s772,s773,s774,s775,s776,s777,s778,s779,s780,s781,s782,s783,s784,s785,s786,s787,s788,s789,s790,s791,s792,p19,p47);
input r827,r828,r829,r830,r831,r832,r833,r834,r835,r836,r837,r838,r839,r840,r841,r842,r843,r844,r845,r846,r847,r848,r849,r850,r851,r852,r853,s737,s738,s739,s740,s741,s742,s743,s744,s745,s746,s747,s748,s749,s750,s751,s752,s753,s754,s755,s756,s757,s758,s759,s760,s761,s762,s763,s764,s765;
output s766,s767,s768,s769,s770,s771,s772,s773,s774,s775,s776,s777,s778,s779,s780,s781,s782,s783,s784,s785,s786,s787,s788,s789,s790,s791,s792,p19,p47;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28;


full_adder fa0(s737,r827,1'b0,p19,d1);
full_adder fa1(s738,r828,d1,s766,d2);
full_adder fa2(s739,r829,d2,s767,d3);
full_adder fa3(s740,r830,d3,s768,d4);
full_adder fa4(s741,r831,d4,s769,d5);
full_adder fa5(s742,r832,d5,s770,d6);
full_adder fa6(s743,r833,d6,s771,d7);
full_adder fa7(s744,r834,d7,s772,d8);
full_adder fa8(s745,r835,d8,s773,d9);
full_adder fa9(s746,r836,d9,s774,d10);
full_adder fa10(s747,r837,d10,s775,d11);
full_adder fa11(s748,r838,d11,s776,d12);
full_adder fa12(s749,r839,d12,s777,d13);
full_adder fa13(s750,r840,d13,s778,d14);
full_adder fa14(s751,r841,d14,s779,d15);
full_adder fa15(s752,r842,d15,s780,d16);
full_adder fa16(s753,r843,d16,s781,d17);
full_adder fa17(s754,r844,d17,s782,d18);
full_adder fa18(s755,r845,d18,s783,d19);
full_adder fa19(s756,r846,d19,s784,d20);
full_adder fa20(s757,r847,d20,s785,d21);
full_adder fa21(s758,r848,d21,s786,d22);
full_adder fa22(s759,r849,d22,s787,d23);
full_adder fa23(s760,r850,d23,s788,d24);
full_adder fa24(s761,r851,d24,s789,d25);
full_adder fa25(s762,r852,d25,s790,d26);
full_adder fa26(s763,r853,d26,s791,d27);
full_adder fa27(s764,1'b0,d27,s792,d28);
full_adder fa28(s765,1'b0,d28,p47,);

endmodule

module stage18(r854,r855,r856,r857,r858,r859,r860,r861,r862,r863,r864,r865,r866,r867,r868,r869,r870,r871,r872,r873,r874,r875,r876,r877,r878,s766,s767,s768,s769,s770,s771,s772,s773,s774,s775,s776,s777,s778,s779,s780,s781,s782,s783,s784,s785,s786,s787,s788,s789,s790,s791,s792,s793,s794,s795,s796,s797,s798,s799,s800,s801,s802,s803,s804,s805,s806,s807,s808,s809,s810,s811,s812,s813,s814,s815,s816,s817,p20,p46);
input r854,r855,r856,r857,r858,r859,r860,r861,r862,r863,r864,r865,r866,r867,r868,r869,r870,r871,r872,r873,r874,r875,r876,r877,r878,s766,s767,s768,s769,s770,s771,s772,s773,s774,s775,s776,s777,s778,s779,s780,s781,s782,s783,s784,s785,s786,s787,s788,s789,s790,s791,s792;
output s793,s794,s795,s796,s797,s798,s799,s800,s801,s802,s803,s804,s805,s806,s807,s808,s809,s810,s811,s812,s813,s814,s815,s816,s817,p20,p46;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26;


full_adder fa0(s766,r854,1'b0,p20,d1);
full_adder fa1(s767,r855,d1,s793,d2);
full_adder fa2(s768,r856,d2,s794,d3);
full_adder fa3(s769,r857,d3,s795,d4);
full_adder fa4(s770,r858,d4,s796,d5);
full_adder fa5(s771,r859,d5,s797,d6);
full_adder fa6(s772,r860,d6,s798,d7);
full_adder fa7(s773,r861,d7,s799,d8);
full_adder fa8(s774,r862,d8,s800,d9);
full_adder fa9(s775,r863,d9,s801,d10);
full_adder fa10(s776,r864,d10,s802,d11);
full_adder fa11(s777,r865,d11,s803,d12);
full_adder fa12(s778,r866,d12,s804,d13);
full_adder fa13(s779,r867,d13,s805,d14);
full_adder fa14(s780,r868,d14,s806,d15);
full_adder fa15(s781,r869,d15,s807,d16);
full_adder fa16(s782,r870,d16,s808,d17);
full_adder fa17(s783,r871,d17,s809,d18);
full_adder fa18(s784,r872,d18,s810,d19);
full_adder fa19(s785,r873,d19,s811,d20);
full_adder fa20(s786,r874,d20,s812,d21);
full_adder fa21(s787,r875,d21,s813,d22);
full_adder fa22(s788,r876,d22,s814,d23);
full_adder fa23(s789,r877,d23,s815,d24);
full_adder fa24(s790,r878,d24,s816,d25);
full_adder fa25(s791,1'b0,d25,s817,d26);
full_adder fa26(s792,1'b0,d26,p46,);

endmodule

module stage19(r879,r880,r881,r882,r883,r884,r885,r886,r887,r888,r889,r890,r891,r892,r893,r894,r895,r896,r897,r898,r899,r900,r901,s793,s794,s795,s796,s797,s798,s799,s800,s801,s802,s803,s804,s805,s806,s807,s808,s809,s810,s811,s812,s813,s814,s815,s816,s817,s818,s819,s820,s821,s822,s823,s824,s825,s826,s827,s828,s829,s830,s831,s832,s833,s834,s835,s836,s837,s838,s839,s840,p21,p45);
input r879,r880,r881,r882,r883,r884,r885,r886,r887,r888,r889,r890,r891,r892,r893,r894,r895,r896,r897,r898,r899,r900,r901,s793,s794,s795,s796,s797,s798,s799,s800,s801,s802,s803,s804,s805,s806,s807,s808,s809,s810,s811,s812,s813,s814,s815,s816,s817;
output s818,s819,s820,s821,s822,s823,s824,s825,s826,s827,s828,s829,s830,s831,s832,s833,s834,s835,s836,s837,s838,s839,s840,p21,p45;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24;


full_adder fa0(s793,r879,1'b0,p21,d1);
full_adder fa1(s794,r880,d1,s818,d2);
full_adder fa2(s795,r881,d2,s819,d3);
full_adder fa3(s796,r882,d3,s820,d4);
full_adder fa4(s797,r883,d4,s821,d5);
full_adder fa5(s798,r884,d5,s822,d6);
full_adder fa6(s799,r885,d6,s823,d7);
full_adder fa7(s800,r886,d7,s824,d8);
full_adder fa8(s801,r887,d8,s825,d9);
full_adder fa9(s802,r888,d9,s826,d10);
full_adder fa10(s803,r889,d10,s827,d11);
full_adder fa11(s804,r890,d11,s828,d12);
full_adder fa12(s805,r891,d12,s829,d13);
full_adder fa13(s806,r892,d13,s830,d14);
full_adder fa14(s807,r893,d14,s831,d15);
full_adder fa15(s808,r894,d15,s832,d16);
full_adder fa16(s809,r895,d16,s833,d17);
full_adder fa17(s810,r896,d17,s834,d18);
full_adder fa18(s811,r897,d18,s835,d19);
full_adder fa19(s812,r898,d19,s836,d20);
full_adder fa20(s813,r899,d20,s837,d21);
full_adder fa21(s814,r900,d21,s838,d22);
full_adder fa22(s815,r901,d22,s839,d23);
full_adder fa23(s816,1'b0,d23,s840,d24);
full_adder fa24(s817,1'b0,d24,p45,);

endmodule

module stage20(r902,r903,r904,r905,r906,r907,r908,r909,r910,r911,r912,r913,r914,r915,r916,r917,r918,r919,r920,r921,r922,s818,s819,s820,s821,s822,s823,s824,s825,s826,s827,s828,s829,s830,s831,s832,s833,s834,s835,s836,s837,s838,s839,s840,s841,s842,s843,s844,s845,s846,s847,s848,s849,s850,s851,s852,s853,s854,s855,s856,s857,s858,s859,s860,s861,p22,p44);
input r902,r903,r904,r905,r906,r907,r908,r909,r910,r911,r912,r913,r914,r915,r916,r917,r918,r919,r920,r921,r922,s818,s819,s820,s821,s822,s823,s824,s825,s826,s827,s828,s829,s830,s831,s832,s833,s834,s835,s836,s837,s838,s839,s840;
output s841,s842,s843,s844,s845,s846,s847,s848,s849,s850,s851,s852,s853,s854,s855,s856,s857,s858,s859,s860,s861,p22,p44;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22;


full_adder fa0(s818,r902,1'b0,p22,d1);
full_adder fa1(s819,r903,d1,s841,d2);
full_adder fa2(s820,r904,d2,s842,d3);
full_adder fa3(s821,r905,d3,s843,d4);
full_adder fa4(s822,r906,d4,s844,d5);
full_adder fa5(s823,r907,d5,s845,d6);
full_adder fa6(s824,r908,d6,s846,d7);
full_adder fa7(s825,r909,d7,s847,d8);
full_adder fa8(s826,r910,d8,s848,d9);
full_adder fa9(s827,r911,d9,s849,d10);
full_adder fa10(s828,r912,d10,s850,d11);
full_adder fa11(s829,r913,d11,s851,d12);
full_adder fa12(s830,r914,d12,s852,d13);
full_adder fa13(s831,r915,d13,s853,d14);
full_adder fa14(s832,r916,d14,s854,d15);
full_adder fa15(s833,r917,d15,s855,d16);
full_adder fa16(s834,r918,d16,s856,d17);
full_adder fa17(s835,r919,d17,s857,d18);
full_adder fa18(s836,r920,d18,s858,d19);
full_adder fa19(s837,r921,d19,s859,d20);
full_adder fa20(s838,r922,d20,s860,d21);
full_adder fa21(s839,1'b0,d21,s861,d22);
full_adder fa22(s840,1'b0,d22,p44,);

endmodule

module stage21(r923,r924,r925,r926,r927,r928,r929,r930,r931,r932,r933,r934,r935,r936,r937,r938,r939,r940,r941,s841,s842,s843,s844,s845,s846,s847,s848,s849,s850,s851,s852,s853,s854,s855,s856,s857,s858,s859,s860,s861,s862,s863,s864,s865,s866,s867,s868,s869,s870,s871,s872,s873,s874,s875,s876,s877,s878,s879,s880,p23,p43);
input r923,r924,r925,r926,r927,r928,r929,r930,r931,r932,r933,r934,r935,r936,r937,r938,r939,r940,r941,s841,s842,s843,s844,s845,s846,s847,s848,s849,s850,s851,s852,s853,s854,s855,s856,s857,s858,s859,s860,s861;
output s862,s863,s864,s865,s866,s867,s868,s869,s870,s871,s872,s873,s874,s875,s876,s877,s878,s879,s880,p23,p43;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20;


full_adder fa0(s841,r923,1'b0,p23,d1);
full_adder fa1(s842,r924,d1,s862,d2);
full_adder fa2(s843,r925,d2,s863,d3);
full_adder fa3(s844,r926,d3,s864,d4);
full_adder fa4(s845,r927,d4,s865,d5);
full_adder fa5(s846,r928,d5,s866,d6);
full_adder fa6(s847,r929,d6,s867,d7);
full_adder fa7(s848,r930,d7,s868,d8);
full_adder fa8(s849,r931,d8,s869,d9);
full_adder fa9(s850,r932,d9,s870,d10);
full_adder fa10(s851,r933,d10,s871,d11);
full_adder fa11(s852,r934,d11,s872,d12);
full_adder fa12(s853,r935,d12,s873,d13);
full_adder fa13(s854,r936,d13,s874,d14);
full_adder fa14(s855,r937,d14,s875,d15);
full_adder fa15(s856,r938,d15,s876,d16);
full_adder fa16(s857,r939,d16,s877,d17);
full_adder fa17(s858,r940,d17,s878,d18);
full_adder fa18(s859,r941,d18,s879,d19);
full_adder fa19(s860,1'b0,d19,s880,d20);
full_adder fa20(s861,1'b0,d20,p43,);

endmodule

module stage22(r942,r943,r944,r945,r946,r947,r948,r949,r950,r951,r952,r953,r954,r955,r956,r957,r958,s862,s863,s864,s865,s866,s867,s868,s869,s870,s871,s872,s873,s874,s875,s876,s877,s878,s879,s880,s881,s882,s883,s884,s885,s886,s887,s888,s889,s890,s891,s892,s893,s894,s895,s896,s897,p24,p42);
input r942,r943,r944,r945,r946,r947,r948,r949,r950,r951,r952,r953,r954,r955,r956,r957,r958,s862,s863,s864,s865,s866,s867,s868,s869,s870,s871,s872,s873,s874,s875,s876,s877,s878,s879,s880;
output s881,s882,s883,s884,s885,s886,s887,s888,s889,s890,s891,s892,s893,s894,s895,s896,s897,p24,p42;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18;


full_adder fa0(s862,r942,1'b0,p24,d1);
full_adder fa1(s863,r943,d1,s881,d2);
full_adder fa2(s864,r944,d2,s882,d3);
full_adder fa3(s865,r945,d3,s883,d4);
full_adder fa4(s866,r946,d4,s884,d5);
full_adder fa5(s867,r947,d5,s885,d6);
full_adder fa6(s868,r948,d6,s886,d7);
full_adder fa7(s869,r949,d7,s887,d8);
full_adder fa8(s870,r950,d8,s888,d9);
full_adder fa9(s871,r951,d9,s889,d10);
full_adder fa10(s872,r952,d10,s890,d11);
full_adder fa11(s873,r953,d11,s891,d12);
full_adder fa12(s874,r954,d12,s892,d13);
full_adder fa13(s875,r955,d13,s893,d14);
full_adder fa14(s876,r956,d14,s894,d15);
full_adder fa15(s877,r957,d15,s895,d16);
full_adder fa16(s878,r958,d16,s896,d17);
full_adder fa17(s879,1'b0,d17,s897,d18);
full_adder fa18(s880,1'b0,d18,p42,);

endmodule

module stage23(r959,r960,r961,r962,r963,r964,r965,r966,r967,r968,r969,r970,r971,r972,r973,s881,s882,s883,s884,s885,s886,s887,s888,s889,s890,s891,s892,s893,s894,s895,s896,s897,s898,s899,s900,s901,s902,s903,s904,s905,s906,s907,s908,s909,s910,s911,s912,p25,p41);
input r959,r960,r961,r962,r963,r964,r965,r966,r967,r968,r969,r970,r971,r972,r973,s881,s882,s883,s884,s885,s886,s887,s888,s889,s890,s891,s892,s893,s894,s895,s896,s897;
output s898,s899,s900,s901,s902,s903,s904,s905,s906,s907,s908,s909,s910,s911,s912,p25,p41;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16;


full_adder fa0(s881,r959,1'b0,p25,d1);
full_adder fa1(s882,r960,d1,s898,d2);
full_adder fa2(s883,r961,d2,s899,d3);
full_adder fa3(s884,r962,d3,s900,d4);
full_adder fa4(s885,r963,d4,s901,d5);
full_adder fa5(s886,r964,d5,s902,d6);
full_adder fa6(s887,r965,d6,s903,d7);
full_adder fa7(s888,r966,d7,s904,d8);
full_adder fa8(s889,r967,d8,s905,d9);
full_adder fa9(s890,r968,d9,s906,d10);
full_adder fa10(s891,r969,d10,s907,d11);
full_adder fa11(s892,r970,d11,s908,d12);
full_adder fa12(s893,r971,d12,s909,d13);
full_adder fa13(s894,r972,d13,s910,d14);
full_adder fa14(s895,r973,d14,s911,d15);
full_adder fa15(s896,1'b0,d15,s912,d16);
full_adder fa16(s897,1'b0,d16,p41,);

endmodule

module stage24(r974,r975,r976,r977,r978,r979,r980,r981,r982,r983,r984,r985,r986,s898,s899,s900,s901,s902,s903,s904,s905,s906,s907,s908,s909,s910,s911,s912,s913,s914,s915,s916,s917,s918,s919,s920,s921,s922,s923,s924,s925,p26,p40);
input r974,r975,r976,r977,r978,r979,r980,r981,r982,r983,r984,r985,r986,s898,s899,s900,s901,s902,s903,s904,s905,s906,s907,s908,s909,s910,s911,s912;
output s913,s914,s915,s916,s917,s918,s919,s920,s921,s922,s923,s924,s925,p26,p40;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14;


full_adder fa0(s898,r974,1'b0,p26,d1);
full_adder fa1(s899,r975,d1,s913,d2);
full_adder fa2(s900,r976,d2,s914,d3);
full_adder fa3(s901,r977,d3,s915,d4);
full_adder fa4(s902,r978,d4,s916,d5);
full_adder fa5(s903,r979,d5,s917,d6);
full_adder fa6(s904,r980,d6,s918,d7);
full_adder fa7(s905,r981,d7,s919,d8);
full_adder fa8(s906,r982,d8,s920,d9);
full_adder fa9(s907,r983,d9,s921,d10);
full_adder fa10(s908,r984,d10,s922,d11);
full_adder fa11(s909,r985,d11,s923,d12);
full_adder fa12(s910,r986,d12,s924,d13);
full_adder fa13(s911,1'b0,d13,s925,d14);
full_adder fa14(s912,1'b0,d14,p40,);

endmodule

module stage25(r987,r988,r989,r990,r991,r992,r993,r994,r995,r996,r997,s913,s914,s915,s916,s917,s918,s919,s920,s921,s922,s923,s924,s925,s926,s927,s928,s929,s930,s931,s932,s933,s934,s935,s936,p27,p39);
input r987,r988,r989,r990,r991,r992,r993,r994,r995,r996,r997,s913,s914,s915,s916,s917,s918,s919,s920,s921,s922,s923,s924,s925;
output s926,s927,s928,s929,s930,s931,s932,s933,s934,s935,s936,p27,p39;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12;


full_adder fa0(s913,r987,1'b0,p27,d1);
full_adder fa1(s914,r988,d1,s926,d2);
full_adder fa2(s915,r989,d2,s927,d3);
full_adder fa3(s916,r990,d3,s928,d4);
full_adder fa4(s917,r991,d4,s929,d5);
full_adder fa5(s918,r992,d5,s930,d6);
full_adder fa6(s919,r993,d6,s931,d7);
full_adder fa7(s920,r994,d7,s932,d8);
full_adder fa8(s921,r995,d8,s933,d9);
full_adder fa9(s922,r996,d9,s934,d10);
full_adder fa10(s923,r997,d10,s935,d11);
full_adder fa11(s924,1'b0,d11,s936,d12);
full_adder fa12(s925,1'b0,d12,p39,);

endmodule

module stage26(r998,r999,r1000,r1001,r1002,r1003,r1004,r1005,r1006,s926,s927,s928,s929,s930,s931,s932,s933,s934,s935,s936,s937,s938,s939,s940,s941,s942,s943,s944,s945,p28,p38);
input r998,r999,r1000,r1001,r1002,r1003,r1004,r1005,r1006,s926,s927,s928,s929,s930,s931,s932,s933,s934,s935,s936;
output s937,s938,s939,s940,s941,s942,s943,s944,s945,p28,p38;
wire d1,d2,d3,d4,d5,d6,d7,d8,d9,d10;


full_adder fa0(s926,r998,1'b0,p28,d1);
full_adder fa1(s927,r999,d1,s937,d2);
full_adder fa2(s928,r1000,d2,s938,d3);
full_adder fa3(s929,r1001,d3,s939,d4);
full_adder fa4(s930,r1002,d4,s940,d5);
full_adder fa5(s931,r1003,d5,s941,d6);
full_adder fa6(s932,r1004,d6,s942,d7);
full_adder fa7(s933,r1005,d7,s943,d8);
full_adder fa8(s934,r1006,d8,s944,d9);
full_adder fa9(s935,1'b0,d9,s945,d10);
full_adder fa10(s936,1'b0,d10,p38,);

endmodule

module stage27(r1007,r1008,r1009,r1010,r1011,r1012,r1013,s937,s938,s939,s940,s941,s942,s943,s944,s945,s946,s947,s948,s949,s950,s951,s952,p29,p37);
input r1007,r1008,r1009,r1010,r1011,r1012,r1013,s937,s938,s939,s940,s941,s942,s943,s944,s945;
output s946,s947,s948,s949,s950,s951,s952,p29,p37;
wire d1,d2,d3,d4,d5,d6,d7,d8;


full_adder fa0(s937,r1007,1'b0,p29,d1);
full_adder fa1(s938,r1008,d1,s946,d2);
full_adder fa2(s939,r1009,d2,s947,d3);
full_adder fa3(s940,r1010,d3,s948,d4);
full_adder fa4(s941,r1011,d4,s949,d5);
full_adder fa5(s942,r1012,d5,s950,d6);
full_adder fa6(s943,r1013,d6,s951,d7);
full_adder fa7(s944,1'b0,d7,s952,d8);
full_adder fa8(s945,1'b0,d8,p37,);

endmodule

module stage28(r1014,r1015,r1016,r1017,r1018,s946,s947,s948,s949,s950,s951,s952,s953,s954,s955,s956,s957,p30,p36);
input r1014,r1015,r1016,r1017,r1018,s946,s947,s948,s949,s950,s951,s952;
output s953,s954,s955,s956,s957,p30,p36;
wire d1,d2,d3,d4,d5,d6;


full_adder fa0(s946,r1014,1'b0,p30,d1);
full_adder fa1(s947,r1015,d1,s953,d2);
full_adder fa2(s948,r1016,d2,s954,d3);
full_adder fa3(s949,r1017,d3,s955,d4);
full_adder fa4(s950,r1018,d4,s956,d5);
full_adder fa5(s951,1'b0,d5,s957,d6);
full_adder fa6(s952,1'b0,d6,p36,);

endmodule

module stage29(r1019,r1020,r1021,s953,s954,s955,s956,s957,s958,s959,s960,p31,p35);
input r1019,r1020,r1021,s953,s954,s955,s956,s957;
output s958,s959,s960,p31,p35;
wire d1,d2,d3,d4;


full_adder fa0(s953,r1019,1'b0,p31,d1);
full_adder fa1(s954,r1020,d1,s958,d2);
full_adder fa2(s955,r1021,d2,s959,d3);
full_adder fa3(s956,1'b0,d3,s960,d4);
full_adder fa4(s957,1'b0,d4,p35,);

endmodule

module stage30(r1022,s958,s959,s960,p32,p33,p34);
input r1022,s958,s959,s960;
output p32,p33,p34;
wire d1,d2;


full_adder fa0(s958,r1022,1'b0,p32,d1);
full_adder fa1(s959,1'b0,d1,p33,d2);
full_adder fa2(s960,1'b0,d2,p34,);

endmodule
