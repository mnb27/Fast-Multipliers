`timescale 1ns / 1ps

module FinalSum(p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,ans);
input p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64;
output reg [63:0]ans;

always@(*)begin
ans[0] <= p1;
ans[1] <= p2;
ans[2] <= p3;
ans[3] <= p4;
ans[4] <= p5;
ans[5] <= p6;
ans[6] <= p7;
ans[7] <= p8;
ans[8] <= p9;
ans[9] <= p10;
ans[10] <= p11;
ans[11] <= p12;
ans[12] <= p13;
ans[13] <= p14;
ans[14] <= p15;
ans[15] <= p16;
ans[16] <= p17;
ans[17] <= p18;
ans[18] <= p19;
ans[19] <= p20;
ans[20] <= p21;
ans[21] <= p22;
ans[22] <= p23;
ans[23] <= p24;
ans[24] <= p25;
ans[25] <= p26;
ans[26] <= p27;
ans[27] <= p28;
ans[28] <= p29;
ans[29] <= p30;
ans[30] <= p31;
ans[31] <= p32;
ans[32] <= p33;
ans[33] <= p34;
ans[34] <= p35;
ans[35] <= p36;
ans[36] <= p37;
ans[37] <= p38;
ans[38] <= p39;
ans[39] <= p40;
ans[40] <= p41;
ans[41] <= p42;
ans[42] <= p43;
ans[43] <= p44;
ans[44] <= p45;
ans[45] <= p46;
ans[46] <= p47;
ans[47] <= p48;
ans[48] <= p49;
ans[49] <= p50;
ans[50] <= p51;
ans[51] <= p52;
ans[52] <= p53;
ans[53] <= p54;
ans[54] <= p55;
ans[55] <= p56;
ans[56] <= p57;
ans[57] <= p58;
ans[58] <= p59;
ans[59] <= p60;
ans[60] <= p61;
ans[61] <= p62;
ans[62] <= p63;
ans[63] <= p64;

end

endmodule
